VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

UNITS
  DATABASE MICRONS 2000 ;
END UNITS

PROPERTYDEFINITIONS
    LAYER LEF58_CORNERSPACING STRING ;
END PROPERTYDEFINITIONS

CLEARANCEMEASURE EUCLIDEAN ;
MANUFACTURINGGRID 0.0005 ;
USEMINSPACING OBS ON ;

LAYER Metal1
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.10 0.10 ;
  WIDTH 0.05 ;
  AREA 0.0115 ;
  MINWIDTH 0.05 ;
  SPACINGTABLE
    PARALLELRUNLENGTH  0.0 0.22 0.47 0.63 1.50
    WIDTH 0.0         0.05 0.05 0.05 0.05 0.05
    WIDTH 0.10        0.05 0.06 0.06 0.06 0.06
    WIDTH 0.28        0.05 0.10 0.10 0.10 0.10
    WIDTH 0.47        0.05 0.10 0.13 0.13 0.13
    WIDTH 0.63        0.05 0.10 0.13 0.15 0.15
    WIDTH 1.50        0.05 0.10 0.13 0.15 0.50 ;
  SPACING 0.06 ENDOFLINE 0.06 WITHIN 0.025 ;
END Metal1

LAYER Via1
  TYPE CUT ;
  SPACING 0.075 ;
  WIDTH 0.05 ;
END Via1

LAYER Metal2
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.10 0.10 ;
  WIDTH 0.05 ;
  AREA 0.014 ;
  MINWIDTH 0.05 ;
  SPACINGTABLE
    PARALLELRUNLENGTH  0.0 0.22 0.47 0.63 1.5
    WIDTH 0.0         0.05 0.05 0.05 0.05 0.05
    WIDTH 0.09        0.05 0.06 0.06 0.06 0.06
    WIDTH 0.16        0.05 0.10 0.10 0.10 0.10
    WIDTH 0.47        0.05 0.10 0.13 0.13 0.13
    WIDTH 0.63        0.05 0.10 0.13 0.15 0.15
    WIDTH 1.5         0.05 0.10 0.13 0.15 0.50 ;
  SPACING 0.08 ENDOFLINE 0.08 WITHIN 0.025 ;
  SPACING 0.10 ENDOFLINE 0.08 WITHIN 0.025 PARALLELEDGE 0.10 WITHIN 0.025 ;
  PROPERTY LEF58_CORNERSPACING "CORNERSPACING CONVEXCORNER EXCEPTEOL 0.08
    WIDTH 0.00 SPACING 0.10
    WIDTH 0.20 SPACING 0.20
    WIDTH 0.50 SPACING 0.30 ;" ;
END Metal2

LAYER Via2
  TYPE CUT ;
  SPACING 0.075 ;
  WIDTH 0.05 ;
  SPACING 0.155 ADJACENTCUTS 3 WITHIN 0.200 ;
END Via2

LAYER Metal3
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.10 0.10 ;
  WIDTH 0.05 ;
  AREA 0.017 ;
  MINWIDTH 0.05 ;
  SPACINGTABLE
    PARALLELRUNLENGTH  0.0 0.22 0.47 0.63 1.5
    WIDTH 0.0         0.05 0.05 0.05 0.05 0.05
    WIDTH 0.09        0.05 0.06 0.06 0.06 0.06
    WIDTH 0.16        0.05 0.10 0.10 0.10 0.10
    WIDTH 0.47        0.05 0.10 0.13 0.13 0.13
    WIDTH 0.63        0.05 0.10 0.13 0.15 0.15
    WIDTH 1.5         0.05 0.10 0.13 0.15 0.50 ;
  SPACING 0.08 ENDOFLINE 0.08 WITHIN 0.025 ;
  SPACING 0.10 ENDOFLINE 0.08 WITHIN 0.025 PARALLELEDGE 0.10 WITHIN 0.025 ;
  PROPERTY LEF58_CORNERSPACING "CORNERSPACING CONVEXCORNER EXCEPTEOL 0.08
    WIDTH 0.00 SPACING 0.10
    WIDTH 0.20 SPACING 0.20
    WIDTH 0.50 SPACING 0.30 ;" ;
END Metal3

LAYER Via3
  TYPE CUT ;
  SPACING 0.075 ;
  WIDTH 0.05 ;
  SPACING 0.155 ADJACENTCUTS 3 WITHIN 0.200 ;
END Via3

LAYER Metal4
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.10 0.10 ;
  WIDTH 0.05 ;
  AREA 0.017 ;
  MINWIDTH 0.05 ;
  SPACINGTABLE
    PARALLELRUNLENGTH  0.0 0.22 0.47 0.63 1.5
    WIDTH 0.0         0.05 0.05 0.05 0.05 0.05
    WIDTH 0.09        0.05 0.06 0.06 0.06 0.06
    WIDTH 0.16        0.05 0.10 0.10 0.10 0.10
    WIDTH 0.47        0.05 0.10 0.13 0.13 0.13
    WIDTH 0.63        0.05 0.10 0.13 0.15 0.15
    WIDTH 1.5         0.05 0.10 0.13 0.15 0.50 ;
  SPACING 0.08 ENDOFLINE 0.08 WITHIN 0.025 ;
  SPACING 0.10 ENDOFLINE 0.08 WITHIN 0.025 PARALLELEDGE 0.10 WITHIN 0.025 ;
  PROPERTY LEF58_CORNERSPACING "CORNERSPACING CONVEXCORNER EXCEPTEOL 0.08
    WIDTH 0.00 SPACING 0.10
    WIDTH 0.20 SPACING 0.20
    WIDTH 0.50 SPACING 0.30 ;" ;
END Metal4

LAYER Via4
  TYPE CUT ;
  SPACING 0.075 ;
  WIDTH 0.05 ;
  SPACING 0.155 ADJACENTCUTS 3 WITHIN 0.200 ;
END Via4

LAYER Metal5
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.10 0.10 ;
  WIDTH 0.05 ;
  AREA 0.017 ;
  MINWIDTH 0.05 ;
  SPACINGTABLE
    PARALLELRUNLENGTH  0.0 0.22 0.47 0.63 1.5
    WIDTH 0.0         0.05 0.05 0.05 0.05 0.05
    WIDTH 0.09        0.05 0.06 0.06 0.06 0.06
    WIDTH 0.16        0.05 0.10 0.10 0.10 0.10
    WIDTH 0.47        0.05 0.10 0.13 0.13 0.13
    WIDTH 0.63        0.05 0.10 0.13 0.15 0.15
    WIDTH 1.5         0.05 0.10 0.13 0.15 0.50 ;
  SPACING 0.08 ENDOFLINE 0.08 WITHIN 0.025 ;
  SPACING 0.10 ENDOFLINE 0.08 WITHIN 0.025 PARALLELEDGE 0.10 WITHIN 0.025 ;
  PROPERTY LEF58_CORNERSPACING "CORNERSPACING CONVEXCORNER EXCEPTEOL 0.08
    WIDTH 0.00 SPACING 0.10
    WIDTH 0.20 SPACING 0.20
    WIDTH 0.50 SPACING 0.30 ;" ;
END Metal5

LAYER Via5
  TYPE CUT ;
  SPACING 0.075 ;
  WIDTH 0.05 ;
  SPACING 0.155 ADJACENTCUTS 3 WITHIN 0.200 ;
END Via5

LAYER Metal6
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.15 0.15 ;
  WIDTH 0.07 ;
  AREA 0.025 ;
  MINWIDTH 0.07 ;
  SPACINGTABLE
    PARALLELRUNLENGTH  0.0 0.22 0.47 0.63 1.5
    WIDTH 0.0         0.08 0.08 0.08 0.08 0.08
    WIDTH 0.10        0.08 0.12 0.12 0.12 0.12
    WIDTH 0.16        0.08 0.12 0.15 0.15 0.15
    WIDTH 0.47        0.08 0.12 0.15 0.18 0.18
    WIDTH 0.63        0.08 0.12 0.15 0.18 0.25
    WIDTH 1.5         0.08 0.12 0.15 0.18 0.50 ;
  SPACING 0.10 ENDOFLINE 0.10 WITHIN 0.035 ;
  SPACING 0.12 ENDOFLINE 0.10 WITHIN 0.035 PARALLELEDGE 0.12 WITHIN 0.035 ;
  PROPERTY LEF58_CORNERSPACING "CORNERSPACING CONVEXCORNER EXCEPTEOL 0.08
    WIDTH 0.00 SPACING 0.10
    WIDTH 0.20 SPACING 0.20
    WIDTH 0.50 SPACING 0.30 ;" ;
END Metal6

LAYER Via6
  TYPE CUT ;
  SPACING 0.10 ;
  WIDTH 0.07 ;
  SPACING 0.20 ADJACENTCUTS 3 WITHIN 0.25 ;
END Via6

LAYER Metal7
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.15 0.15 ;
  WIDTH 0.07 ;
  AREA 0.025 ;
  MINWIDTH 0.07 ;
  SPACINGTABLE
    PARALLELRUNLENGTH  0.0 0.22 0.47 0.63 1.5
    WIDTH 0.0         0.08 0.08 0.08 0.08 0.08
    WIDTH 0.10        0.08 0.12 0.12 0.12 0.12
    WIDTH 0.16        0.08 0.12 0.15 0.15 0.15
    WIDTH 0.47        0.08 0.12 0.15 0.18 0.18
    WIDTH 0.63        0.08 0.12 0.15 0.18 0.25
    WIDTH 1.5         0.08 0.12 0.15 0.18 0.50 ;
  SPACING 0.10 ENDOFLINE 0.10 WITHIN 0.035 ;
  SPACING 0.12 ENDOFLINE 0.10 WITHIN 0.035 PARALLELEDGE 0.12 WITHIN 0.035 ;
  PROPERTY LEF58_CORNERSPACING "CORNERSPACING CONVEXCORNER EXCEPTEOL 0.08
    WIDTH 0.00 SPACING 0.10
    WIDTH 0.20 SPACING 0.20
    WIDTH 0.50 SPACING 0.30 ;" ;
END Metal7

LAYER Via7
  TYPE CUT ;
  SPACING 0.10 ;
  WIDTH 0.07 ;
  SPACING 0.20 ADJACENTCUTS 3 WITHIN 0.25 ;
END Via7

LAYER Metal8
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.2 0.2 ;
  WIDTH 0.10 ;
  AREA 0.052 ;
  MINWIDTH 0.10 ;
  SPACINGTABLE
    PARALLELRUNLENGTH 0.0 0.22 0.47 0.63 1.5
    WIDTH 0	     0.10 0.10 0.10 0.10 0.10
    WIDTH 0.2	     0.10 0.15 0.15 0.15 0.15
    WIDTH 0.4	     0.10 0.15 0.20 0.20 0.20
    WIDTH 1.5	     0.10 0.15 0.20 0.30 0.50 ;
  SPACING 0.12 ENDOFLINE 0.12 WITHIN 0.035 ;
END Metal8

LAYER Via8
  TYPE CUT ;
  SPACING 0.15 ;
  WIDTH 0.10 ;
END Via8

LAYER Metal9
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.2 0.2 ;
  WIDTH 0.10 ;
  AREA 0.052 ;
  MINWIDTH 0.10 ;
  SPACINGTABLE
    PARALLELRUNLENGTH 0.0 0.22 0.47 0.63 1.5
    WIDTH 0	     0.10 0.10 0.10 0.10 0.10
    WIDTH 0.2	     0.10 0.15 0.15 0.15 0.15
    WIDTH 0.4	     0.10 0.15 0.20 0.20 0.20
    WIDTH 1.5	     0.10 0.15 0.20 0.30 0.50 ;
  SPACING 0.12 ENDOFLINE 0.12 WITHIN 0.035 ;
END Metal9

LAYER OVERLAP
  TYPE OVERLAP ;
END OVERLAP

VIA VIA12_1C DEFAULT 
    LAYER Metal1 ;
        RECT -0.025000 -0.055000 0.025000 0.055000 ;
    LAYER Via1 ;
        RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal2 ;
        RECT -0.055000 -0.025000 0.055000 0.025000 ;
END VIA12_1C

VIA VIA12_1C_H DEFAULT 
    LAYER Metal1 ;
        RECT -0.055000 -0.025000 0.055000 0.025000 ;
    LAYER Via1 ;
        RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal2 ;
        RECT -0.055000 -0.025000 0.055000 0.025000 ;
END VIA12_1C_H

VIA VIA12_1C_V DEFAULT 
    LAYER Metal1 ;
        RECT -0.025000 -0.055000 0.025000 0.055000 ;
    LAYER Via1 ;
        RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal2 ;
        RECT -0.025000 -0.055000 0.025000 0.055000 ;
END VIA12_1C_V

VIA VIA12_PG
    LAYER Metal1 ;
        RECT -0.350000 -0.050000 0.350000 0.050000 ;
    LAYER Via1 ;
        RECT -0.325000 -0.025000 -0.275000 0.025000 ;
        RECT -0.175000 -0.025000 -0.125000 0.025000 ;
        RECT -0.025000 -0.025000 0.025000 0.025000 ;
        RECT 0.125000 -0.025000 0.175000 0.025000 ;
        RECT 0.275000 -0.025000 0.325000 0.025000 ;
    LAYER Metal2 ;
        RECT -0.350000 -0.050000 0.350000 0.050000 ;
END VIA12_PG

VIA VIA23_1C DEFAULT 
    LAYER Metal2 ;
        RECT -0.055000 -0.025000 0.055000 0.025000 ;
    LAYER Via2 ;
        RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal3 ;
        RECT -0.025000 -0.055000 0.025000 0.055000 ;
END VIA23_1C

VIA VIA23_1C_H DEFAULT 
    LAYER Metal2 ;
        RECT -0.055000 -0.025000 0.055000 0.025000 ;
    LAYER Via2 ;
        RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal3 ;
        RECT -0.055000 -0.025000 0.055000 0.025000 ;
END VIA23_1C_H

VIA VIA23_1C_V DEFAULT 
    LAYER Metal2 ;
        RECT -0.025000 -0.055000 0.025000 0.055000 ;
    LAYER Via2 ;
        RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal3 ;
        RECT -0.025000 -0.055000 0.025000 0.055000 ;
END VIA23_1C_V

VIA VIA23_1ST_E DEFAULT 
    LAYER Metal2 ;
        RECT -0.055000 -0.025000 0.325000 0.025000 ;
    LAYER Via2 ;
        RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal3 ;
        RECT -0.025000 -0.055000 0.025000 0.055000 ;
END VIA23_1ST_E

VIA VIA23_1ST_W DEFAULT 
    LAYER Metal2 ;
        RECT -0.325000 -0.025000 0.055000 0.025000 ;
    LAYER Via2 ;
        RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal3 ;
        RECT -0.025000 -0.055000 0.025000 0.055000 ;
END VIA23_1ST_W

VIA VIA23_PG
    LAYER Metal2 ;
        RECT -0.350000 -0.050000 0.350000 0.050000 ;
    LAYER Via2 ;
        RECT -0.325000 -0.025000 -0.275000 0.025000 ;
        RECT -0.175000 -0.025000 -0.125000 0.025000 ;
        RECT -0.025000 -0.025000 0.025000 0.025000 ;
        RECT 0.125000 -0.025000 0.175000 0.025000 ;
        RECT 0.275000 -0.025000 0.325000 0.025000 ;
    LAYER Metal3 ;
        RECT -0.350000 -0.050000 0.350000 0.050000 ;
END VIA23_PG

VIA VIA34_1C DEFAULT 
    LAYER Metal3 ;
        RECT -0.025000 -0.055000 0.025000 0.055000 ;
    LAYER Via3 ;
        RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal4 ;
        RECT -0.055000 -0.025000 0.055000 0.025000 ;
END VIA34_1C

VIA VIA34_1C_H DEFAULT 
    LAYER Metal3 ;
        RECT -0.055000 -0.025000 0.055000 0.025000 ;
    LAYER Via3 ;
        RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal4 ;
        RECT -0.055000 -0.025000 0.055000 0.025000 ;
END VIA34_1C_H

VIA VIA34_1C_V DEFAULT 
    LAYER Metal3 ;
        RECT -0.025000 -0.055000 0.025000 0.055000 ;
    LAYER Via3 ;
        RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal4 ;
        RECT -0.025000 -0.055000 0.025000 0.055000 ;
END VIA34_1C_V

VIA VIA34_1ST_N DEFAULT 
    LAYER Metal3 ;
        RECT -0.025000 -0.055000 0.025000 0.325000 ;
    LAYER Via3 ;
        RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal4 ;
        RECT -0.055000 -0.025000 0.055000 0.025000 ;
END VIA34_1ST_N

VIA VIA34_1ST_S DEFAULT 
    LAYER Metal3 ;
        RECT -0.025000 -0.325000 0.025000 0.055000 ;
    LAYER Via3 ;
        RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal4 ;
        RECT -0.055000 -0.025000 0.055000 0.025000 ;
END VIA34_1ST_S

VIA VIA34_PG
    LAYER Metal3 ;
        RECT -0.350000 -0.050000 0.350000 0.050000 ;
    LAYER Via3 ;
        RECT -0.325000 -0.025000 -0.275000 0.025000 ;
        RECT -0.175000 -0.025000 -0.125000 0.025000 ;
        RECT -0.025000 -0.025000 0.025000 0.025000 ;
        RECT 0.125000 -0.025000 0.175000 0.025000 ;
        RECT 0.275000 -0.025000 0.325000 0.025000 ;
    LAYER Metal4 ;
        RECT -0.350000 -0.050000 0.350000 0.050000 ;
END VIA34_PG

VIA VIA45_1C DEFAULT 
    LAYER Metal4 ;
        RECT -0.055000 -0.025000 0.055000 0.025000 ;
    LAYER Via4 ;
        RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal5 ;
        RECT -0.025000 -0.055000 0.025000 0.055000 ;
END VIA45_1C

VIA VIA45_PG
    LAYER Metal4 ;
        RECT -0.200000 -0.050000 0.200000 0.050000 ;
    LAYER Via4 ;
        RECT -0.175000 -0.025000 -0.125000 0.025000 ;
        RECT -0.025000 -0.025000 0.025000 0.025000 ;
        RECT 0.125000 -0.025000 0.175000 0.025000 ;
    LAYER Metal5 ;
        RECT -0.200000 -0.050000 0.200000 0.050000 ;
END VIA45_PG

VIA VIA5_0_VH DEFAULT 
    LAYER Metal5 ;
        RECT -0.035000 -0.065000 0.035000 0.065000 ;
    LAYER Via5 ;
        RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal6 ;
        RECT -0.065000 -0.035000 0.065000 0.035000 ;
END VIA5_0_VH

VIA VIA56_PG
    LAYER Metal5 ;
        RECT -0.150000 -0.150000 0.150000 0.150000 ;
    LAYER Via5 ;
        RECT -0.150000 -0.150000 -0.100000 -0.100000 ;
        RECT -0.150000 0.100000 -0.100000 0.150000 ;
        RECT 0.100000 0.100000 0.150000 0.150000 ;
        RECT 0.100000 -0.150000 0.150000 -0.100000 ;
    LAYER Metal6 ;
        RECT -0.150000 -0.150000 0.150000 0.150000 ;
END VIA56_PG

VIA VIA6_0_HV DEFAULT 
    LAYER Metal6 ;
        RECT -0.065000 -0.035000 0.065000 0.035000 ;
    LAYER Via6 ;
        RECT -0.035000 -0.035000 0.035000 0.035000 ;
    LAYER Metal7 ;
        RECT -0.035000 -0.065000 0.035000 0.065000 ;
END VIA6_0_HV

VIA VIA67_PG
    LAYER Metal6 ;
        RECT -0.170000 -0.170000 0.170000 0.170000 ;
    LAYER Via6 ;
        RECT -0.170000 -0.170000 -0.100000 -0.100000 ;
        RECT -0.170000 0.100000 -0.100000 0.170000 ;
        RECT 0.100000 0.100000 0.170000 0.170000 ;
        RECT 0.100000 -0.170000 0.170000 -0.100000 ;
    LAYER Metal7 ;
        RECT -0.170000 -0.170000 0.170000 0.170000 ;
END VIA67_PG

VIA VIA7_0_VH DEFAULT 
    LAYER Metal7 ;
        RECT -0.050000 -0.260000 0.050000 0.260000 ;
    LAYER Via7 ;
        RECT -0.050000 -0.050000 0.050000 0.050000 ;
    LAYER Metal8 ;
        RECT -0.260000 -0.050000 0.260000 0.050000 ;
END VIA7_0_VH

VIA VIA78_PG
    LAYER Metal7 ;
        RECT -0.170000 -0.170000 0.170000 0.170000 ;
    LAYER Via7 ;
        RECT -0.170000 -0.170000 -0.100000 -0.100000 ;
        RECT -0.170000 0.100000 -0.100000 0.170000 ;
        RECT 0.100000 0.100000 0.170000 0.170000 ;
        RECT 0.100000 -0.170000 0.170000 -0.100000 ;
    LAYER Metal8 ;
        RECT -0.170000 -0.170000 0.170000 0.170000 ;
END VIA78_PG

VIA VIA8_0_HV DEFAULT 
    LAYER Metal8 ;
        RECT -0.260000 -0.050000 0.260000 0.050000 ;
    LAYER Via8 ;
        RECT -0.050000 -0.050000 0.050000 0.050000 ;
    LAYER Metal9 ;
        RECT -0.050000 -0.260000 0.050000 0.260000 ;
END VIA8_0_HV

VIA VIA12_2C_W DEFAULT
    LAYER Metal1 ;
	RECT -0.150000 -0.055000 0.025000 0.055000 ;
    LAYER Via1 ;
	RECT -0.025000 -0.025000 0.025000 0.025000 ;
	RECT -0.150000 -0.025000 -0.100000 0.025000 ;
    LAYER Metal2 ;
	RECT -0.180000 -0.025000 0.055000 0.025000 ;
END VIA12_2C_W

VIA VIA12_2C_CH DEFAULT
    LAYER Metal1 ;
	RECT -0.087500 -0.055000 0.087500 0.055000 ;
    LAYER Via1 ;
	RECT 0.037500 -0.025000 0.087500 0.025000 ;
	RECT -0.087500 -0.025000 -0.037500 0.025000 ;
    LAYER Metal2 ;
	RECT -0.117500 -0.025000 0.117500 0.025000 ;
END VIA12_2C_CH

VIA VIA12_2C_E DEFAULT
    LAYER Metal1 ;
	RECT -0.025000 -0.055000 0.150000 0.055000 ;
    LAYER Via1 ;
	RECT 0.100000 -0.025000 0.150000 0.025000 ;
	RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal2 ;
	RECT -0.055000 -0.025000 0.180000 0.025000 ;
END VIA12_2C_E

VIA VIA12_2C_S DEFAULT
    LAYER Metal1 ;
	RECT -0.025000 -0.180000 0.025000 0.055000 ;
    LAYER Via1 ;
	RECT -0.025000 -0.025000 0.025000 0.025000 ;
	RECT -0.025000 -0.150000 0.025000 -0.100000 ;
    LAYER Metal2 ;
	RECT -0.055000 -0.150000 0.055000 0.025000 ;
END VIA12_2C_S

VIA VIA12_2C_CV DEFAULT
    LAYER Metal1 ;
	RECT -0.025000 -0.117500 0.025000 0.117500 ;
    LAYER Via1 ;
	RECT -0.025000 0.037500 0.025000 0.087500 ;
	RECT -0.025000 -0.087500 0.025000 -0.037500 ;
    LAYER Metal2 ;
	RECT -0.055000 -0.087500 0.055000 0.087500 ;
END VIA12_2C_CV

VIA VIA12_2C_N DEFAULT
    LAYER Metal1 ;
	RECT -0.025000 -0.055000 0.025000 0.180000 ;
    LAYER Via1 ;
	RECT -0.025000 0.100000 0.025000 0.150000 ;
	RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal2 ;
	RECT -0.055000 -0.025000 0.055000 0.150000 ;
END VIA12_2C_N

VIA VIA23_2C_W DEFAULT
    LAYER Metal2 ;
	RECT -0.180000 -0.025000 0.055000 0.025000 ;
    LAYER Via2 ;
	RECT -0.025000 -0.025000 0.025000 0.025000 ;
	RECT -0.150000 -0.025000 -0.100000 0.025000 ;
    LAYER Metal3 ;
	RECT -0.150000 -0.055000 0.025000 0.055000 ;
END VIA23_2C_W

VIA VIA23_2C_CH DEFAULT
    LAYER Metal2 ;
	RECT -0.117500 -0.025000 0.117500 0.025000 ;
    LAYER Via2 ;
	RECT 0.037500 -0.025000 0.087500 0.025000 ;
	RECT -0.087500 -0.025000 -0.037500 0.025000 ;
    LAYER Metal3 ;
	RECT -0.087500 -0.055000 0.087500 0.055000 ;
END VIA23_2C_CH

VIA VIA23_2C_E DEFAULT
    LAYER Metal2 ;
	RECT -0.055000 -0.025000 0.180000 0.025000 ;
    LAYER Via2 ;
	RECT 0.100000 -0.025000 0.150000 0.025000 ;
	RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal3 ;
	RECT -0.025000 -0.055000 0.150000 0.055000 ;
END VIA23_2C_E

VIA VIA23_2C_S DEFAULT
    LAYER Metal2 ;
	RECT -0.055000 -0.150000 0.055000 0.025000 ;
    LAYER Via2 ;
	RECT -0.025000 -0.025000 0.025000 0.025000 ;
	RECT -0.025000 -0.150000 0.025000 -0.100000 ;
    LAYER Metal3 ;
	RECT -0.025000 -0.180000 0.025000 0.055000 ;
END VIA23_2C_S

VIA VIA23_2C_CV DEFAULT
    LAYER Metal2 ;
	RECT -0.055000 -0.087500 0.055000 0.087500 ;
    LAYER Via2 ;
	RECT -0.025000 0.037500 0.025000 0.087500 ;
	RECT -0.025000 -0.087500 0.025000 -0.037500 ;
    LAYER Metal3 ;
	RECT -0.025000 -0.117500 0.025000 0.117500 ;
END VIA23_2C_CV

VIA VIA23_2C_N DEFAULT
    LAYER Metal2 ;
	RECT -0.055000 -0.025000 0.055000 0.150000 ;
    LAYER Via2 ;
	RECT -0.025000 0.100000 0.025000 0.150000 ;
	RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal3 ;
	RECT -0.025000 -0.055000 0.025000 0.180000 ;
END VIA23_2C_N

VIA VIA34_2C_W DEFAULT
    LAYER Metal3 ;
	RECT -0.150000 -0.055000 0.025000 0.055000 ;
    LAYER Via3 ;
	RECT -0.025000 -0.025000 0.025000 0.025000 ;
	RECT -0.150000 -0.025000 -0.100000 0.025000 ;
    LAYER Metal4 ;
	RECT -0.180000 -0.025000 0.055000 0.025000 ;
END VIA34_2C_W

VIA VIA34_2C_CH DEFAULT
    LAYER Metal3 ;
	RECT -0.087500 -0.055000 0.087500 0.055000 ;
    LAYER Via3 ;
	RECT 0.037500 -0.025000 0.087500 0.025000 ;
	RECT -0.087500 -0.025000 -0.037500 0.025000 ;
    LAYER Metal4 ;
	RECT -0.117500 -0.025000 0.117500 0.025000 ;
END VIA34_2C_CH

VIA VIA34_2C_E DEFAULT
    LAYER Metal3 ;
	RECT -0.025000 -0.055000 0.150000 0.055000 ;
    LAYER Via3 ;
	RECT 0.100000 -0.025000 0.150000 0.025000 ;
	RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal4 ;
	RECT -0.055000 -0.025000 0.180000 0.025000 ;
END VIA34_2C_E

VIA VIA34_2C_S DEFAULT
    LAYER Metal3 ;
	RECT -0.025000 -0.180000 0.025000 0.055000 ;
    LAYER Via3 ;
	RECT -0.025000 -0.025000 0.025000 0.025000 ;
	RECT -0.025000 -0.150000 0.025000 -0.100000 ;
    LAYER Metal4 ;
	RECT -0.055000 -0.150000 0.055000 0.025000 ;
END VIA34_2C_S

VIA VIA34_2C_CV DEFAULT
    LAYER Metal3 ;
	RECT -0.025000 -0.117500 0.025000 0.117500 ;
    LAYER Via3 ;
	RECT -0.025000 0.037500 0.025000 0.087500 ;
	RECT -0.025000 -0.087500 0.025000 -0.037500 ;
    LAYER Metal4 ;
	RECT -0.055000 -0.087500 0.055000 0.087500 ;
END VIA34_2C_CV

VIA VIA34_2C_N DEFAULT
    LAYER Metal3 ;
	RECT -0.025000 -0.055000 0.025000 0.180000 ;
    LAYER Via3 ;
	RECT -0.025000 0.100000 0.025000 0.150000 ;
	RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal4 ;
	RECT -0.055000 -0.025000 0.055000 0.150000 ;
END VIA34_2C_N

VIA VIA45_2C_W DEFAULT
    LAYER Metal4 ;
	RECT -0.180000 -0.025000 0.055000 0.025000 ;
    LAYER Via4 ;
	RECT -0.025000 -0.025000 0.025000 0.025000 ;
	RECT -0.150000 -0.025000 -0.100000 0.025000 ;
    LAYER Metal5 ;
	RECT -0.150000 -0.055000 0.025000 0.055000 ;
END VIA45_2C_W

VIA VIA45_2C_CH DEFAULT
    LAYER Metal4 ;
	RECT -0.117500 -0.025000 0.117500 0.025000 ;
    LAYER Via4 ;
	RECT 0.037500 -0.025000 0.087500 0.025000 ;
	RECT -0.087500 -0.025000 -0.037500 0.025000 ;
    LAYER Metal5 ;
	RECT -0.087500 -0.055000 0.087500 0.055000 ;
END VIA45_2C_CH

VIA VIA45_2C_E DEFAULT
    LAYER Metal4 ;
	RECT -0.055000 -0.025000 0.180000 0.025000 ;
    LAYER Via4 ;
	RECT 0.100000 -0.025000 0.150000 0.025000 ;
	RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal5 ;
	RECT -0.025000 -0.055000 0.150000 0.055000 ;
END VIA45_2C_E

VIA VIA45_2C_S DEFAULT
    LAYER Metal4 ;
	RECT -0.055000 -0.150000 0.055000 0.025000 ;
    LAYER Via4 ;
	RECT -0.025000 -0.025000 0.025000 0.025000 ;
	RECT -0.025000 -0.150000 0.025000 -0.100000 ;
    LAYER Metal5 ;
	RECT -0.025000 -0.180000 0.025000 0.055000 ;
END VIA45_2C_S

VIA VIA45_2C_CV DEFAULT
    LAYER Metal4 ;
	RECT -0.055000 -0.087500 0.055000 0.087500 ;
    LAYER Via4 ;
	RECT -0.025000 0.037500 0.025000 0.087500 ;
	RECT -0.025000 -0.087500 0.025000 -0.037500 ;
    LAYER Metal5 ;
	RECT -0.025000 -0.117500 0.025000 0.117500 ;
END VIA45_2C_CV

VIA VIA45_2C_N DEFAULT
    LAYER Metal4 ;
	RECT -0.055000 -0.025000 0.055000 0.150000 ;
    LAYER Via4 ;
	RECT -0.025000 0.100000 0.025000 0.150000 ;
	RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal5 ;
	RECT -0.025000 -0.055000 0.025000 0.180000 ;
END VIA45_2C_N

VIA VIA56_2C_W DEFAULT
    LAYER Metal5 ;
	RECT -0.150000 -0.055000 0.025000 0.055000 ;
    LAYER Via5 ;
	RECT -0.025000 -0.025000 0.025000 0.025000 ;
	RECT -0.150000 -0.025000 -0.100000 0.025000 ;
    LAYER Metal6 ;
	RECT -0.180000 -0.025000 0.055000 0.025000 ;
END VIA56_2C_W

VIA VIA56_2C_CH DEFAULT
    LAYER Metal5 ;
	RECT -0.087500 -0.055000 0.087500 0.055000 ;
    LAYER Via5 ;
	RECT 0.037500 -0.025000 0.087500 0.025000 ;
	RECT -0.087500 -0.025000 -0.037500 0.025000 ;
    LAYER Metal6 ;
	RECT -0.117500 -0.025000 0.117500 0.025000 ;
END VIA56_2C_CH

VIA VIA56_2C_E DEFAULT
    LAYER Metal5 ;
	RECT -0.025000 -0.055000 0.150000 0.055000 ;
    LAYER Via5 ;
	RECT 0.100000 -0.025000 0.150000 0.025000 ;
	RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal6 ;
	RECT -0.055000 -0.025000 0.180000 0.025000 ;
END VIA56_2C_E

VIA VIA56_2C_S DEFAULT
    LAYER Metal5 ;
	RECT -0.025000 -0.180000 0.025000 0.055000 ;
    LAYER Via5 ;
	RECT -0.025000 -0.025000 0.025000 0.025000 ;
	RECT -0.025000 -0.150000 0.025000 -0.100000 ;
    LAYER Metal6 ;
	RECT -0.055000 -0.150000 0.055000 0.025000 ;
END VIA56_2C_S

VIA VIA56_2C_CV DEFAULT
    LAYER Metal5 ;
	RECT -0.025000 -0.117500 0.025000 0.117500 ;
    LAYER Via5 ;
	RECT -0.025000 0.037500 0.025000 0.087500 ;
	RECT -0.025000 -0.087500 0.025000 -0.037500 ;
    LAYER Metal6 ;
	RECT -0.055000 -0.087500 0.055000 0.087500 ;
END VIA56_2C_CV

VIA VIA56_2C_N DEFAULT
    LAYER Metal5 ;
	RECT -0.025000 -0.055000 0.025000 0.180000 ;
    LAYER Via5 ;
	RECT -0.025000 0.100000 0.025000 0.150000 ;
	RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal6 ;
	RECT -0.055000 -0.025000 0.055000 0.150000 ;
END VIA56_2C_N

VIA VIA67_2C_W DEFAULT
    LAYER Metal6 ;
	RECT -0.235000 -0.035000 0.065000 0.035000 ;
    LAYER Via6 ;
	RECT -0.035000 -0.035000 0.035000 0.035000 ;
	RECT -0.205000 -0.035000 -0.135000 0.035000 ;
    LAYER Metal7 ;
	RECT -0.205000 -0.065000 0.035000 0.065000 ;
END VIA67_2C_W

VIA VIA67_2C_CH DEFAULT
    LAYER Metal6 ;
	RECT -0.150000 -0.035000 0.150000 0.035000 ;
    LAYER Via6 ;
	RECT 0.050000 -0.035000 0.120000 0.035000 ;
	RECT -0.120000 -0.035000 -0.050000 0.035000 ;
    LAYER Metal7 ;
	RECT -0.120000 -0.065000 0.120000 0.065000 ;
END VIA67_2C_CH

VIA VIA67_2C_E DEFAULT
    LAYER Metal6 ;
	RECT -0.065000 -0.035000 0.235000 0.035000 ;
    LAYER Via6 ;
	RECT 0.135000 -0.035000 0.205000 0.035000 ;
	RECT -0.035000 -0.035000 0.035000 0.035000 ;
    LAYER Metal7 ;
	RECT -0.035000 -0.065000 0.205000 0.065000 ;
END VIA67_2C_E

VIA VIA67_2C_S DEFAULT
    LAYER Metal6 ;
	RECT -0.065000 -0.205000 0.065000 0.035000 ;
    LAYER Via6 ;
	RECT -0.035000 -0.035000 0.035000 0.035000 ;
	RECT -0.035000 -0.205000 0.035000 -0.135000 ;
    LAYER Metal7 ;
	RECT -0.035000 -0.235000 0.035000 0.065000 ;
END VIA67_2C_S

VIA VIA67_2C_CV DEFAULT
    LAYER Metal6 ;
	RECT -0.065000 -0.120000 0.065000 0.120000 ;
    LAYER Via6 ;
	RECT -0.035000 0.050000 0.035000 0.120000 ;
	RECT -0.035000 -0.120000 0.035000 -0.050000 ;
    LAYER Metal7 ;
	RECT -0.035000 -0.150000 0.035000 0.150000 ;
END VIA67_2C_CV

VIA VIA67_2C_N DEFAULT
    LAYER Metal6 ;
	RECT -0.065000 -0.035000 0.065000 0.205000 ;
    LAYER Via6 ;
	RECT -0.035000 0.135000 0.035000 0.205000 ;
	RECT -0.035000 -0.035000 0.035000 0.035000 ;
    LAYER Metal7 ;
	RECT -0.035000 -0.065000 0.035000 0.235000 ;
END VIA67_2C_N

VIA VIA78_2C_W DEFAULT
    LAYER Metal7 ;
	RECT -0.205000 -0.065000 0.035000 0.065000 ;
    LAYER Via7 ;
	RECT -0.035000 -0.035000 0.035000 0.035000 ;
	RECT -0.205000 -0.035000 -0.135000 0.035000 ;
    LAYER Metal8 ;
	RECT -0.235000 -0.035000 0.065000 0.035000 ;
END VIA78_2C_W

VIA VIA78_2C_CH DEFAULT
    LAYER Metal7 ;
	RECT -0.120000 -0.065000 0.120000 0.065000 ;
    LAYER Via7 ;
	RECT 0.050000 -0.035000 0.120000 0.035000 ;
	RECT -0.120000 -0.035000 -0.050000 0.035000 ;
    LAYER Metal8 ;
	RECT -0.150000 -0.035000 0.150000 0.035000 ;
END VIA78_2C_CH

VIA VIA78_2C_E DEFAULT
    LAYER Metal7 ;
	RECT -0.035000 -0.065000 0.205000 0.065000 ;
    LAYER Via7 ;
	RECT 0.135000 -0.035000 0.205000 0.035000 ;
	RECT -0.035000 -0.035000 0.035000 0.035000 ;
    LAYER Metal8 ;
	RECT -0.065000 -0.035000 0.235000 0.035000 ;
END VIA78_2C_E

VIA VIA78_2C_S DEFAULT
    LAYER Metal7 ;
	RECT -0.035000 -0.235000 0.035000 0.065000 ;
    LAYER Via7 ;
	RECT -0.035000 -0.035000 0.035000 0.035000 ;
	RECT -0.035000 -0.205000 0.035000 -0.135000 ;
    LAYER Metal8 ;
	RECT -0.065000 -0.205000 0.065000 0.035000 ;
END VIA78_2C_S

VIA VIA78_2C_CV DEFAULT
    LAYER Metal7 ;
	RECT -0.035000 -0.150000 0.035000 0.150000 ;
    LAYER Via7 ;
	RECT -0.035000 0.050000 0.035000 0.120000 ;
	RECT -0.035000 -0.120000 0.035000 -0.050000 ;
    LAYER Metal8 ;
	RECT -0.065000 -0.120000 0.065000 0.120000 ;
END VIA78_2C_CV

VIA VIA78_2C_N DEFAULT
    LAYER Metal7 ;
	RECT -0.035000 -0.065000 0.035000 0.235000 ;
    LAYER Via7 ;
	RECT -0.035000 0.135000 0.035000 0.205000 ;
	RECT -0.035000 -0.035000 0.035000 0.035000 ;
    LAYER Metal8 ;
	RECT -0.065000 -0.035000 0.065000 0.205000 ;
END VIA78_2C_N

VIARULE M4_M3 GENERATE DEFAULT
  LAYER Metal3 ;
    ENCLOSURE 0.005 0.03 ;
  LAYER Via3 ;
    RECT -0.025 -0.025 0.025 0.025 ;
    SPACING 0.11 BY 0.11 ;
  LAYER Metal4 ;
    ENCLOSURE 0.005 0.03 ;
END M4_M3

VIARULE M5_M4 GENERATE DEFAULT
  LAYER Metal4 ;
    ENCLOSURE 0.005 0.03 ;
  LAYER Via4 ;
    RECT -0.025 -0.025 0.025 0.025 ;
    SPACING 0.11 BY 0.11 ;
  LAYER Metal5 ;
    ENCLOSURE 0.005 0.03 ;
END M5_M4

VIARULE M6_M5 GENERATE DEFAULT
  LAYER Metal5 ;
    ENCLOSURE 0.005 0.03 ;
  LAYER Via5 ;
    RECT -0.025 -0.025 0.025 0.025 ;
    SPACING 0.11 BY 0.11 ;
  LAYER Metal6 ;
    ENCLOSURE 0.005 0.03 ;
END M6_M5

VIARULE M7_M6 GENERATE DEFAULT
  LAYER Metal6 ;
    ENCLOSURE 0.005 0.03 ;
  LAYER Via6 ;
    RECT -0.035 -0.035 0.035 0.035 ;
    SPACING 0.15 BY 0.15 ;
  LAYER Metal7 ;
    ENCLOSURE 0.005 0.03 ;
END M7_M6

VIARULE M8_M7 GENERATE DEFAULT
  LAYER Metal7 ;
    ENCLOSURE 0.005 0.03 ;
  LAYER Via7 ;
    RECT -0.035 -0.035 0.035 0.035 ;
    SPACING 0.15 BY 0.15 ;
  LAYER Metal8 ;
    ENCLOSURE 0.005 0.03 ;
END M8_M7

SITE CoreSite
  CLASS CORE ;
  SIZE 0.1 BY 1.2 ;
END CoreSite


MACRO XOR2X2
    CLASS CORE ;
    FOREIGN XOR2X2 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 1.800000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.574000 0.530000 0.686000 0.630000 ;
        RECT 0.574000 0.454000 0.637000 0.630000 ;
        RECT 0.166000 0.454000 0.229000 0.555000 ;
        RECT 0.869000 0.499000 0.931000 0.585000 ;
        RECT 0.574000 0.530000 0.931000 0.585000 ;
        RECT 0.166000 0.454000 0.637000 0.508000 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.368000 0.564000 0.461000 0.694000 ;
        RECT 0.263000 0.639000 0.326000 0.763000 ;
        RECT 0.239000 0.706000 0.326000 0.763000 ;
        RECT 0.263000 0.639000 0.461000 0.694000 ;
        END
    END B
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 1.800000 1.280000 ;
        RECT 1.437000 1.078000 1.530000 1.280000 ;
        RECT 0.605000 0.905000 0.698000 1.280000 ;
        RECT 0.213000 0.905000 0.305000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 1.800000 0.080000 ;
        RECT 1.440000 -0.080000 1.533000 0.122000 ;
        RECT 0.627000 -0.080000 0.720000 0.122000 ;
        RECT 0.213000 -0.080000 0.305000 0.122000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.655000 0.693000 1.748000 0.998000 ;
        RECT 1.655000 0.171000 1.748000 0.395000 ;
        RECT 1.685000 0.171000 1.748000 0.998000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 0.041000 0.281000 0.142000 0.387000 ;
        RECT 0.818000 0.163000 0.911000 0.261000 ;
        RECT 0.802000 0.717000 0.895000 0.940000 ;
        RECT 1.520000 0.473000 1.621000 0.558000 ;
        RECT 1.015000 0.212000 1.182000 0.293000 ;
        RECT 0.998000 0.783000 1.091000 0.864000 ;
        RECT 0.717000 0.319000 0.810000 0.400000 ;
        RECT 0.420000 0.193000 0.513000 0.274000 ;
        RECT 0.409000 0.824000 0.502000 0.905000 ;
        RECT 0.041000 0.950000 0.138000 1.031000 ;
        RECT 0.041000 0.683000 0.142000 0.764000 ;
        RECT 1.520000 0.212000 1.583000 0.558000 ;
        RECT 1.376000 0.520000 1.439000 0.994000 ;
        RECT 1.245000 0.336000 1.308000 0.802000 ;
        RECT 0.994000 0.368000 1.057000 0.708000 ;
        RECT 0.832000 0.654000 0.895000 0.994000 ;
        RECT 0.439000 0.765000 0.502000 0.905000 ;
        RECT 0.041000 0.281000 0.104000 1.031000 ;
        RECT 1.120000 0.212000 1.182000 0.838000 ;
        RECT 0.884000 0.206000 0.946000 0.423000 ;
        RECT 1.015000 0.212000 1.583000 0.267000 ;
        RECT 0.998000 0.783000 1.182000 0.838000 ;
        RECT 0.884000 0.368000 1.057000 0.423000 ;
        RECT 0.832000 0.939000 1.439000 0.994000 ;
        RECT 0.717000 0.206000 0.946000 0.261000 ;
        RECT 0.439000 0.765000 0.895000 0.820000 ;
        RECT 0.420000 0.206000 0.832000 0.261000 ;
        RECT 0.138000 0.332000 0.810000 0.387000 ;
        RECT 0.041000 0.332000 0.513000 0.387000 ;
        RECT 0.832000 0.654000 1.057000 0.708000 ;
        RECT 0.884000 0.163000 0.911000 0.423000 ;
    END
END XOR2X2

MACRO XNOR2X2
    CLASS CORE ;
    FOREIGN XNOR2X2 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 2.000000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.059000 0.468000 1.123000 0.585000 ;
        RECT 0.811000 0.530000 0.875000 0.630000 ;
        RECT 0.584000 0.454000 0.647000 0.630000 ;
        RECT 0.168000 0.454000 0.231000 0.555000 ;
        RECT 0.584000 0.573000 0.668000 0.630000 ;
        RECT 0.811000 0.530000 1.123000 0.585000 ;
        RECT 0.584000 0.575000 0.875000 0.630000 ;
        RECT 0.168000 0.454000 0.647000 0.508000 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.427000 0.564000 0.521000 0.645000 ;
        RECT 0.402000 0.627000 0.490000 0.694000 ;
        RECT 0.427000 0.564000 0.490000 0.694000 ;
        RECT 0.266000 0.639000 0.329000 0.763000 ;
        RECT 0.241000 0.706000 0.329000 0.763000 ;
        RECT 0.266000 0.639000 0.490000 0.694000 ;
        END
    END B
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 2.000000 1.280000 ;
        RECT 0.694000 0.905000 0.788000 1.280000 ;
        RECT 1.634000 1.078000 1.727000 1.280000 ;
        RECT 0.287000 0.905000 0.380000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 2.000000 0.080000 ;
        RECT 1.647000 -0.080000 1.741000 0.122000 ;
        RECT 0.716000 -0.080000 0.810000 0.122000 ;
        RECT 0.292000 -0.080000 0.386000 0.122000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.854000 0.693000 1.948000 0.998000 ;
        RECT 1.857000 0.171000 1.950000 0.395000 ;
        RECT 1.884000 0.171000 1.948000 0.998000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 1.207000 0.196000 1.376000 0.302000 ;
        RECT 0.927000 0.717000 1.022000 0.940000 ;
        RECT 0.041000 0.281000 0.143000 0.376000 ;
        RECT 1.718000 0.471000 1.820000 0.558000 ;
        RECT 1.190000 0.783000 1.284000 0.864000 ;
        RECT 0.862000 0.308000 0.956000 0.389000 ;
        RECT 0.507000 0.186000 0.601000 0.267000 ;
        RECT 0.496000 0.824000 0.590000 0.905000 ;
        RECT 0.041000 0.950000 0.139000 1.031000 ;
        RECT 0.041000 0.683000 0.143000 0.764000 ;
        RECT 1.439000 0.306000 1.503000 0.802000 ;
        RECT 1.023000 0.199000 1.087000 0.412000 ;
        RECT 0.526000 0.765000 0.590000 0.905000 ;
        RECT 0.041000 0.281000 0.105000 1.031000 ;
        RECT 1.718000 0.196000 1.781000 0.558000 ;
        RECT 1.572000 0.520000 1.635000 0.994000 ;
        RECT 1.313000 0.196000 1.376000 0.838000 ;
        RECT 1.186000 0.357000 1.249000 0.708000 ;
        RECT 0.959000 0.654000 1.022000 0.994000 ;
        RECT 1.207000 0.196000 1.781000 0.251000 ;
        RECT 1.190000 0.783000 1.376000 0.838000 ;
        RECT 1.023000 0.357000 1.249000 0.412000 ;
        RECT 0.959000 0.939000 1.635000 0.994000 ;
        RECT 0.862000 0.199000 1.087000 0.254000 ;
        RECT 0.601000 0.199000 1.023000 0.254000 ;
        RECT 0.526000 0.765000 1.022000 0.820000 ;
        RECT 0.507000 0.199000 1.022000 0.254000 ;
        RECT 0.139000 0.321000 0.956000 0.376000 ;
        RECT 0.041000 0.321000 0.601000 0.376000 ;
        RECT 0.959000 0.654000 1.249000 0.708000 ;
    END
END XNOR2X2

MACRO SEDFFTRX2
    CLASS CORE ;
    FOREIGN SEDFFTRX2 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 7.000000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER Metal1 ;
        RECT 3.208000 0.439000 3.443000 0.494000 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.457000 0.439000 1.624000 0.524000 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 2.128000 0.433000 2.241000 0.550000 ;
        END
    END E
    PIN Q
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 6.821000 0.346000 6.920000 0.427000 ;
        RECT 6.810000 0.656000 6.901000 0.737000 ;
        RECT 6.810000 0.656000 6.920000 0.724000 ;
        RECT 6.859000 0.306000 6.920000 0.724000 ;
        RECT 6.859000 0.306000 6.943000 0.361000 ;
        RECT 6.859000 0.306000 6.901000 0.737000 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 6.482000 0.346000 6.572000 0.427000 ;
        RECT 6.471000 0.656000 6.561000 0.737000 ;
        RECT 6.496000 0.346000 6.572000 0.439000 ;
        RECT 6.496000 0.573000 6.561000 0.737000 ;
        RECT 6.496000 0.346000 6.557000 0.737000 ;
        RECT 6.496000 0.573000 6.593000 0.627000 ;
        END
    END QN
    PIN RN
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.212000 0.356000 0.293000 0.494000 ;
        RECT 0.170000 0.343000 0.260000 0.424000 ;
        RECT 0.170000 0.356000 0.293000 0.424000 ;
        RECT 0.212000 0.343000 0.260000 0.494000 ;
        END
    END RN
    PIN SE
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.379000 0.514000 0.488000 0.633000 ;
        END
    END SE
    PIN SI
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.697000 0.150000 0.838000 0.258000 ;
        END
    END SI
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 4.164000 1.078000 4.413000 1.280000 ;
        RECT 0.000000 1.120000 7.000000 1.280000 ;
        RECT 5.841000 0.863000 5.953000 1.280000 ;
        RECT 6.641000 0.971000 6.731000 1.280000 ;
        RECT 4.897000 1.078000 4.987000 1.280000 ;
        RECT 3.281000 1.008000 3.371000 1.280000 ;
        RECT 2.227000 1.008000 2.317000 1.280000 ;
        RECT 1.466000 1.008000 1.556000 1.280000 ;
        RECT 0.398000 1.078000 0.488000 1.280000 ;
        RECT 5.772000 0.863000 6.022000 0.914000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 5.149000 -0.080000 5.398000 0.199000 ;
        RECT 5.144000 -0.080000 5.404000 0.118000 ;
        RECT 0.000000 -0.080000 7.000000 0.080000 ;
        RECT 3.648000 -0.080000 3.739000 0.335000 ;
        RECT 0.518000 -0.080000 0.609000 0.197000 ;
        RECT 6.651000 -0.080000 6.741000 0.258000 ;
        RECT 6.052000 -0.080000 6.142000 0.122000 ;
        RECT 4.367000 -0.080000 4.457000 0.274000 ;
        RECT 3.287000 -0.080000 3.377000 0.122000 ;
        RECT 2.255000 -0.080000 2.345000 0.245000 ;
        RECT 1.481000 -0.080000 1.571000 0.122000 ;
        RECT 0.072000 -0.080000 0.162000 0.122000 ;
        END
    END VSS
    OBS
        LAYER Metal1 ;
        RECT 6.153000 0.699000 6.338000 0.887000 ;
        RECT 2.853000 0.645000 2.946000 0.789000 ;
        RECT 6.256000 0.162000 6.346000 0.386000 ;
        RECT 6.153000 0.699000 6.243000 0.952000 ;
        RECT 0.048000 0.874000 0.138000 0.994000 ;
        RECT 2.483000 0.456000 2.585000 0.543000 ;
        RECT 1.144000 0.493000 1.322000 0.575000 ;
        RECT 6.126000 0.464000 6.216000 0.545000 ;
        RECT 5.783000 0.419000 5.873000 0.500000 ;
        RECT 5.687000 0.269000 5.778000 0.350000 ;
        RECT 4.770000 0.231000 4.860000 0.312000 ;
        RECT 4.558000 0.221000 4.648000 0.302000 ;
        RECT 4.407000 0.349000 4.497000 0.430000 ;
        RECT 4.184000 0.517000 4.274000 0.598000 ;
        RECT 3.866000 0.301000 3.956000 0.382000 ;
        RECT 3.081000 0.257000 3.171000 0.338000 ;
        RECT 2.846000 0.271000 2.937000 0.352000 ;
        RECT 2.665000 0.645000 2.755000 0.726000 ;
        RECT 2.655000 0.271000 2.746000 0.352000 ;
        RECT 2.469000 0.279000 2.559000 0.360000 ;
        RECT 2.042000 0.293000 2.132000 0.374000 ;
        RECT 1.108000 0.255000 1.198000 0.336000 ;
        RECT 0.732000 0.338000 0.822000 0.419000 ;
        RECT 4.695000 0.379000 4.775000 0.460000 ;
        RECT 4.477000 0.660000 4.619000 0.740000 ;
        RECT 1.294000 0.260000 1.384000 0.340000 ;
        RECT 0.880000 0.657000 0.960000 0.742000 ;
        RECT 6.126000 0.458000 6.202000 0.551000 ;
        RECT 5.783000 0.419000 5.859000 0.506000 ;
        RECT 1.071000 0.693000 1.147000 0.829000 ;
        RECT 4.709000 0.244000 4.775000 0.460000 ;
        RECT 1.259000 0.493000 1.322000 0.694000 ;
        RECT 6.737000 0.505000 6.798000 0.592000 ;
        RECT 6.674000 0.537000 6.735000 0.887000 ;
        RECT 6.277000 0.162000 6.338000 0.887000 ;
        RECT 6.126000 0.282000 6.187000 0.630000 ;
        RECT 5.546000 0.699000 5.607000 0.994000 ;
        RECT 5.424000 0.575000 5.485000 0.817000 ;
        RECT 5.287000 0.451000 5.348000 0.870000 ;
        RECT 5.160000 0.327000 5.221000 0.740000 ;
        RECT 5.038000 0.483000 5.099000 0.746000 ;
        RECT 4.714000 0.244000 4.775000 0.623000 ;
        RECT 4.558000 0.221000 4.619000 0.746000 ;
        RECT 4.215000 0.543000 4.276000 0.727000 ;
        RECT 4.046000 0.192000 4.107000 0.596000 ;
        RECT 3.841000 0.737000 3.902000 0.870000 ;
        RECT 3.801000 0.327000 3.862000 0.485000 ;
        RECT 3.800000 0.542000 3.861000 0.679000 ;
        RECT 3.708000 0.861000 3.769000 0.994000 ;
        RECT 3.678000 0.430000 3.739000 0.792000 ;
        RECT 3.554000 0.735000 3.615000 0.915000 ;
        RECT 3.432000 0.883000 3.493000 1.039000 ;
        RECT 3.041000 0.270000 3.102000 0.665000 ;
        RECT 2.853000 0.271000 2.914000 0.789000 ;
        RECT 2.681000 0.271000 2.742000 0.726000 ;
        RECT 2.665000 0.645000 2.726000 0.789000 ;
        RECT 2.483000 0.279000 2.544000 0.665000 ;
        RECT 1.986000 0.306000 2.047000 0.665000 ;
        RECT 1.861000 0.267000 1.922000 0.789000 ;
        RECT 1.808000 0.640000 1.869000 0.829000 ;
        RECT 1.685000 0.269000 1.746000 0.680000 ;
        RECT 1.261000 0.273000 1.322000 0.694000 ;
        RECT 1.022000 0.281000 1.083000 0.789000 ;
        RECT 0.899000 0.175000 0.960000 0.938000 ;
        RECT 0.732000 0.338000 0.793000 0.725000 ;
        RECT 0.561000 0.939000 0.622000 1.048000 ;
        RECT 0.549000 0.368000 0.610000 0.865000 ;
        RECT 0.374000 0.336000 0.435000 0.423000 ;
        RECT 0.292000 0.161000 0.353000 0.261000 ;
        RECT 0.211000 0.657000 0.272000 0.754000 ;
        RECT 0.048000 0.206000 0.109000 0.994000 ;
        RECT 2.302000 0.468000 2.362000 0.665000 ;
        RECT 4.215000 0.517000 4.274000 0.727000 ;
        RECT 6.674000 0.537000 6.798000 0.592000 ;
        RECT 6.153000 0.832000 6.735000 0.887000 ;
        RECT 5.687000 0.282000 6.187000 0.337000 ;
        RECT 5.546000 0.699000 6.338000 0.754000 ;
        RECT 5.424000 0.575000 6.187000 0.630000 ;
        RECT 5.287000 0.451000 5.859000 0.506000 ;
        RECT 5.160000 0.327000 5.408000 0.382000 ;
        RECT 4.684000 0.568000 4.775000 0.623000 ;
        RECT 4.046000 0.362000 4.497000 0.417000 ;
        RECT 3.841000 0.815000 5.348000 0.870000 ;
        RECT 3.801000 0.327000 3.956000 0.382000 ;
        RECT 3.708000 0.939000 5.607000 0.994000 ;
        RECT 3.678000 0.737000 3.902000 0.792000 ;
        RECT 3.678000 0.430000 3.862000 0.485000 ;
        RECT 2.302000 0.468000 2.421000 0.523000 ;
        RECT 1.656000 0.269000 1.746000 0.324000 ;
        RECT 1.617000 0.625000 1.746000 0.680000 ;
        RECT 1.259000 0.639000 1.355000 0.694000 ;
        RECT 1.071000 0.774000 1.869000 0.829000 ;
        RECT 1.022000 0.281000 1.198000 0.336000 ;
        RECT 0.899000 0.883000 3.493000 0.938000 ;
        RECT 0.899000 0.175000 0.994000 0.230000 ;
        RECT 0.675000 0.670000 0.793000 0.725000 ;
        RECT 0.561000 0.993000 1.364000 1.048000 ;
        RECT 0.374000 0.368000 0.610000 0.423000 ;
        RECT 0.211000 0.699000 0.610000 0.754000 ;
        RECT 0.048000 0.939000 0.622000 0.994000 ;
        RECT 0.048000 0.206000 0.353000 0.261000 ;
        RECT 4.558000 0.692000 5.099000 0.746000 ;
        RECT 4.215000 0.673000 4.619000 0.727000 ;
        RECT 4.004000 0.192000 4.107000 0.246000 ;
        RECT 3.800000 0.542000 4.107000 0.596000 ;
        RECT 3.554000 0.861000 3.769000 0.915000 ;
        RECT 3.432000 0.985000 3.629000 1.039000 ;
        RECT 3.041000 0.611000 3.739000 0.665000 ;
        RECT 2.853000 0.735000 3.615000 0.789000 ;
        RECT 2.427000 0.611000 2.544000 0.665000 ;
        RECT 1.986000 0.611000 2.362000 0.665000 ;
        RECT 1.808000 0.735000 2.726000 0.789000 ;
        RECT 0.549000 0.811000 0.825000 0.865000 ;
        RECT 0.292000 0.161000 0.392000 0.215000 ;
        RECT 2.681000 0.271000 2.726000 0.789000 ;
        RECT 1.294000 0.260000 1.322000 0.694000 ;
        RECT 3.081000 0.257000 3.102000 0.665000 ;
        RECT 1.071000 0.281000 1.083000 0.829000 ;
        RECT 1.861000 0.267000 1.869000 0.829000 ;
        RECT 4.770000 0.231000 4.775000 0.623000 ;
        RECT 2.042000 0.293000 2.047000 0.665000 ;
    END
END SEDFFTRX2

MACRO SEDFFHQX4
    CLASS CORE ;
    FOREIGN SEDFFHQX4 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 6.600000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER Metal1 ;
        RECT 2.421000 0.494000 2.605000 0.575000 ;
        RECT 2.479000 0.494000 2.549000 0.627000 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.079000 0.433000 1.180000 0.564000 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.774000 0.549000 1.874000 0.693000 ;
        RECT 1.704000 0.555000 1.874000 0.610000 ;
        END
    END E
    PIN Q
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 6.246000 0.433000 6.389000 0.733000 ;
        RECT 6.289000 0.433000 6.389000 0.767000 ;
        RECT 6.246000 0.345000 6.336000 0.733000 ;
        RECT 6.289000 0.345000 6.336000 0.767000 ;
        END
    END Q
    PIN SE
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.170000 0.490000 0.291000 0.633000 ;
        END
    END SE
    PIN SI
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.371000 0.167000 0.512000 0.262000 ;
        END
    END SI
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 5.530000 1.078000 5.757000 1.280000 ;
        RECT 2.978000 1.078000 3.220000 1.280000 ;
        RECT 0.000000 1.120000 6.600000 1.280000 ;
        RECT 1.022000 1.078000 1.112000 1.280000 ;
        RECT 0.221000 1.078000 0.311000 1.280000 ;
        RECT 6.428000 1.078000 6.517000 1.280000 ;
        RECT 6.057000 0.735000 6.146000 1.280000 ;
        RECT 2.612000 1.078000 2.701000 1.280000 ;
        RECT 1.729000 1.078000 1.818000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 6.600000 0.080000 ;
        RECT 5.667000 -0.080000 5.757000 0.122000 ;
        RECT 3.343000 -0.080000 3.433000 0.287000 ;
        RECT 2.643000 -0.080000 2.733000 0.122000 ;
        RECT 0.205000 -0.080000 0.295000 0.122000 ;
        RECT 6.425000 -0.080000 6.514000 0.122000 ;
        RECT 6.057000 -0.080000 6.146000 0.364000 ;
        RECT 4.336000 -0.080000 4.425000 0.122000 ;
        RECT 3.936000 -0.080000 4.025000 0.122000 ;
        RECT 1.733000 -0.080000 1.822000 0.122000 ;
        RECT 1.025000 -0.080000 1.114000 0.122000 ;
        END
    END VSS
    OBS
        LAYER Metal1 ;
        RECT 3.684000 0.192000 3.821000 0.355000 ;
        RECT 4.571000 0.301000 4.784000 0.392000 ;
        RECT 5.867000 0.717000 5.957000 0.910000 ;
        RECT 1.958000 0.542000 2.070000 0.631000 ;
        RECT 1.521000 0.526000 1.613000 0.613000 ;
        RECT 0.786000 0.469000 0.886000 0.554000 ;
        RECT 5.687000 0.543000 5.782000 0.627000 ;
        RECT 5.878000 0.507000 6.186000 0.589000 ;
        RECT 2.037000 0.833000 2.126000 0.915000 ;
        RECT 5.867000 0.290000 5.957000 0.371000 ;
        RECT 2.438000 0.231000 2.528000 0.312000 ;
        RECT 0.416000 0.343000 0.505000 0.424000 ;
        RECT 0.395000 0.746000 0.484000 0.827000 ;
        RECT 0.047000 0.343000 0.137000 0.424000 ;
        RECT 2.226000 0.835000 2.316000 0.915000 ;
        RECT 5.867000 0.717000 5.942000 1.007000 ;
        RECT 5.563000 0.301000 5.624000 0.787000 ;
        RECT 5.430000 0.418000 5.491000 0.586000 ;
        RECT 4.671000 0.531000 4.732000 0.898000 ;
        RECT 4.550000 0.692000 4.611000 0.787000 ;
        RECT 4.150000 0.843000 4.211000 0.940000 ;
        RECT 4.150000 0.301000 4.211000 0.787000 ;
        RECT 4.013000 0.508000 4.074000 0.831000 ;
        RECT 3.684000 0.192000 3.745000 0.720000 ;
        RECT 3.547000 0.281000 3.608000 0.831000 ;
        RECT 3.426000 0.357000 3.487000 0.549000 ;
        RECT 3.425000 0.843000 3.486000 0.940000 ;
        RECT 3.250000 0.540000 3.311000 0.682000 ;
        RECT 2.964000 0.844000 3.025000 1.007000 ;
        RECT 2.392000 0.954000 2.453000 1.031000 ;
        RECT 2.268000 0.306000 2.329000 0.899000 ;
        RECT 2.100000 0.687000 2.161000 0.888000 ;
        RECT 1.376000 0.287000 1.437000 0.888000 ;
        RECT 1.242000 0.300000 1.303000 0.725000 ;
        RECT 0.947000 0.202000 1.008000 0.888000 ;
        RECT 0.825000 0.318000 0.886000 0.733000 ;
        RECT 0.609000 0.446000 0.670000 1.008000 ;
        RECT 0.076000 0.746000 0.137000 0.989000 ;
        RECT 0.047000 0.343000 0.108000 0.827000 ;
        RECT 5.878000 0.290000 5.938000 1.007000 ;
        RECT 5.687000 0.192000 5.747000 0.898000 ;
        RECT 4.491000 0.151000 4.551000 0.246000 ;
        RECT 4.278000 0.952000 4.338000 1.050000 ;
        RECT 3.303000 0.952000 3.363000 1.050000 ;
        RECT 3.087000 0.735000 3.147000 0.898000 ;
        RECT 3.033000 0.244000 3.093000 0.680000 ;
        RECT 2.849000 0.257000 2.909000 0.789000 ;
        RECT 2.132000 0.390000 2.192000 0.742000 ;
        RECT 2.079000 0.306000 2.139000 0.445000 ;
        RECT 1.958000 0.150000 2.018000 0.749000 ;
        RECT 1.907000 0.954000 1.967000 1.031000 ;
        RECT 1.832000 0.375000 1.892000 0.482000 ;
        RECT 1.553000 0.302000 1.613000 0.736000 ;
        RECT 1.553000 0.161000 1.613000 0.246000 ;
        RECT 0.829000 0.163000 0.889000 0.257000 ;
        RECT 0.641000 0.343000 0.701000 0.501000 ;
        RECT 0.470000 0.935000 0.530000 1.050000 ;
        RECT 0.416000 0.343000 0.476000 0.827000 ;
        RECT 4.983000 0.732000 5.624000 0.787000 ;
        RECT 4.793000 0.843000 5.747000 0.898000 ;
        RECT 4.625000 0.531000 5.491000 0.586000 ;
        RECT 4.491000 0.151000 4.722000 0.206000 ;
        RECT 4.278000 0.952000 5.942000 1.007000 ;
        RECT 4.150000 0.843000 4.732000 0.898000 ;
        RECT 4.150000 0.732000 4.611000 0.787000 ;
        RECT 4.150000 0.301000 5.624000 0.356000 ;
        RECT 3.684000 0.665000 3.836000 0.720000 ;
        RECT 3.547000 0.776000 4.074000 0.831000 ;
        RECT 3.303000 0.995000 4.338000 1.050000 ;
        RECT 3.250000 0.627000 3.608000 0.682000 ;
        RECT 3.087000 0.843000 3.486000 0.898000 ;
        RECT 3.033000 0.357000 3.487000 0.412000 ;
        RECT 2.986000 0.625000 3.093000 0.680000 ;
        RECT 2.986000 0.244000 3.093000 0.299000 ;
        RECT 2.964000 0.952000 3.363000 1.007000 ;
        RECT 2.849000 0.394000 2.967000 0.449000 ;
        RECT 2.438000 0.257000 2.909000 0.312000 ;
        RECT 2.226000 0.844000 3.025000 0.899000 ;
        RECT 1.958000 0.150000 2.054000 0.205000 ;
        RECT 1.907000 0.976000 2.453000 1.031000 ;
        RECT 1.553000 0.681000 1.657000 0.736000 ;
        RECT 1.553000 0.427000 1.892000 0.482000 ;
        RECT 1.553000 0.302000 1.649000 0.357000 ;
        RECT 1.172000 0.670000 1.303000 0.725000 ;
        RECT 1.172000 0.300000 1.303000 0.355000 ;
        RECT 0.829000 0.202000 1.008000 0.257000 ;
        RECT 0.797000 0.833000 2.161000 0.888000 ;
        RECT 0.797000 0.163000 0.889000 0.218000 ;
        RECT 4.920000 0.192000 5.747000 0.246000 ;
        RECT 3.684000 0.192000 4.551000 0.246000 ;
        RECT 3.425000 0.886000 4.211000 0.940000 ;
        RECT 2.849000 0.735000 3.147000 0.789000 ;
        RECT 2.412000 0.717000 2.909000 0.771000 ;
        RECT 2.392000 0.954000 2.867000 1.008000 ;
        RECT 1.553000 0.192000 2.018000 0.246000 ;
        RECT 1.299000 0.161000 1.613000 0.215000 ;
        RECT 0.609000 0.954000 1.967000 1.008000 ;
        RECT 0.076000 0.935000 0.530000 0.989000 ;
        RECT 2.268000 0.306000 2.316000 0.915000 ;
        RECT 0.076000 0.343000 0.108000 0.989000 ;
        RECT 2.132000 0.390000 2.161000 0.888000 ;
        RECT 0.641000 0.343000 0.670000 1.008000 ;
        RECT 2.100000 0.687000 2.126000 0.915000 ;
        RECT 2.132000 0.306000 2.139000 0.888000 ;
    END
END SEDFFHQX4

MACRO SEDFFHQX2
    CLASS CORE ;
    FOREIGN SEDFFHQX2 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 5.900000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER Metal1 ;
        RECT 2.448000 0.421000 2.628000 0.512000 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.078000 0.433000 1.179000 0.564000 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.772000 0.549000 1.872000 0.693000 ;
        RECT 1.702000 0.555000 1.872000 0.610000 ;
        END
    END E
    PIN Q
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 5.763000 0.652000 5.862000 0.767000 ;
        RECT 5.758000 0.652000 5.863000 0.733000 ;
        RECT 5.758000 0.346000 5.863000 0.427000 ;
        RECT 5.803000 0.346000 5.863000 0.733000 ;
        RECT 5.803000 0.346000 5.862000 0.767000 ;
        END
    END Q
    PIN SE
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.170000 0.490000 0.291000 0.633000 ;
        END
    END SE
    PIN SI
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.371000 0.167000 0.511000 0.262000 ;
        END
    END SI
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 5.900000 1.280000 ;
        RECT 5.579000 1.078000 5.669000 1.280000 ;
        RECT 5.186000 1.078000 5.276000 1.280000 ;
        RECT 1.727000 1.078000 1.817000 1.280000 ;
        RECT 1.021000 1.078000 1.111000 1.280000 ;
        RECT 3.149000 1.078000 3.238000 1.280000 ;
        RECT 0.221000 1.078000 0.310000 1.280000 ;
        RECT 2.624000 0.902000 2.684000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 5.900000 0.080000 ;
        RECT 5.579000 -0.080000 5.669000 0.122000 ;
        RECT 3.340000 -0.080000 3.430000 0.287000 ;
        RECT 1.731000 -0.080000 1.821000 0.122000 ;
        RECT 5.205000 -0.080000 5.294000 0.122000 ;
        RECT 4.311000 -0.080000 4.400000 0.395000 ;
        RECT 3.932000 -0.080000 4.021000 0.342000 ;
        RECT 2.641000 -0.080000 2.730000 0.122000 ;
        RECT 1.024000 -0.080000 1.113000 0.122000 ;
        RECT 0.205000 -0.080000 0.294000 0.122000 ;
        END
    END VSS
    OBS
        LAYER Metal1 ;
        RECT 5.404000 0.748000 5.494000 0.940000 ;
        RECT 1.956000 0.542000 2.068000 0.631000 ;
        RECT 1.520000 0.526000 1.612000 0.613000 ;
        RECT 0.785000 0.469000 0.885000 0.554000 ;
        RECT 5.652000 0.500000 5.741000 0.581000 ;
        RECT 5.404000 0.292000 5.494000 0.373000 ;
        RECT 5.278000 0.543000 5.368000 0.624000 ;
        RECT 4.121000 0.276000 4.211000 0.357000 ;
        RECT 2.983000 0.255000 3.072000 0.336000 ;
        RECT 2.436000 0.231000 2.525000 0.312000 ;
        RECT 1.942000 0.668000 2.031000 0.749000 ;
        RECT 1.566000 0.668000 1.655000 0.749000 ;
        RECT 1.361000 0.287000 1.450000 0.368000 ;
        RECT 1.171000 0.657000 1.261000 0.738000 ;
        RECT 1.171000 0.287000 1.261000 0.368000 ;
        RECT 0.626000 0.343000 0.715000 0.424000 ;
        RECT 0.594000 0.820000 0.684000 0.901000 ;
        RECT 0.455000 0.969000 0.544000 1.050000 ;
        RECT 0.415000 0.343000 0.505000 0.424000 ;
        RECT 0.394000 0.746000 0.484000 0.827000 ;
        RECT 0.047000 0.343000 0.137000 0.424000 ;
        RECT 5.278000 0.543000 5.353000 0.627000 ;
        RECT 4.852000 0.814000 4.927000 0.927000 ;
        RECT 1.956000 0.542000 2.031000 0.749000 ;
        RECT 0.455000 0.935000 0.530000 1.050000 ;
        RECT 2.063000 0.833000 2.190000 0.902000 ;
        RECT 5.432000 0.526000 5.494000 0.940000 ;
        RECT 5.116000 0.683000 5.177000 0.910000 ;
        RECT 5.053000 0.855000 5.114000 1.050000 ;
        RECT 5.031000 0.174000 5.092000 0.268000 ;
        RECT 4.973000 0.573000 5.034000 0.773000 ;
        RECT 4.881000 0.718000 4.942000 0.895000 ;
        RECT 4.840000 0.330000 4.901000 0.649000 ;
        RECT 4.609000 0.261000 4.670000 0.792000 ;
        RECT 4.488000 0.735000 4.549000 0.927000 ;
        RECT 4.472000 0.150000 4.533000 0.242000 ;
        RECT 4.338000 0.594000 4.399000 0.940000 ;
        RECT 3.544000 0.231000 3.605000 0.831000 ;
        RECT 3.030000 0.268000 3.091000 0.650000 ;
        RECT 2.266000 0.306000 2.327000 0.915000 ;
        RECT 2.077000 0.306000 2.138000 0.445000 ;
        RECT 1.956000 0.150000 2.017000 0.749000 ;
        RECT 1.911000 0.954000 1.972000 1.037000 ;
        RECT 1.551000 0.302000 1.612000 0.736000 ;
        RECT 1.551000 0.161000 1.612000 0.246000 ;
        RECT 1.375000 0.287000 1.436000 0.899000 ;
        RECT 0.828000 0.163000 0.889000 0.257000 ;
        RECT 0.824000 0.318000 0.885000 0.733000 ;
        RECT 0.623000 0.820000 0.684000 1.008000 ;
        RECT 0.415000 0.343000 0.476000 0.827000 ;
        RECT 0.076000 0.746000 0.137000 0.989000 ;
        RECT 0.047000 0.343000 0.108000 0.827000 ;
        RECT 5.432000 0.292000 5.492000 0.940000 ;
        RECT 5.105000 0.213000 5.165000 0.627000 ;
        RECT 4.834000 0.150000 4.894000 0.229000 ;
        RECT 4.136000 0.276000 4.196000 0.805000 ;
        RECT 4.010000 0.508000 4.070000 0.831000 ;
        RECT 3.681000 0.289000 3.741000 0.720000 ;
        RECT 3.422000 0.843000 3.482000 0.940000 ;
        RECT 3.418000 0.357000 3.478000 0.462000 ;
        RECT 3.300000 0.954000 3.360000 1.050000 ;
        RECT 2.987000 0.595000 3.047000 0.783000 ;
        RECT 2.866000 0.665000 2.926000 0.898000 ;
        RECT 2.745000 0.776000 2.805000 1.008000 ;
        RECT 2.698000 0.257000 2.758000 0.720000 ;
        RECT 2.130000 0.390000 2.190000 0.902000 ;
        RECT 1.830000 0.375000 1.890000 0.482000 ;
        RECT 1.240000 0.300000 1.300000 0.725000 ;
        RECT 0.947000 0.202000 1.007000 0.899000 ;
        RECT 0.626000 0.343000 0.686000 0.501000 ;
        RECT 0.609000 0.446000 0.669000 0.901000 ;
        RECT 5.432000 0.526000 5.741000 0.581000 ;
        RECT 5.053000 0.855000 5.494000 0.910000 ;
        RECT 5.031000 0.213000 5.165000 0.268000 ;
        RECT 4.881000 0.718000 5.034000 0.773000 ;
        RECT 4.840000 0.330000 5.038000 0.385000 ;
        RECT 4.834000 0.174000 5.092000 0.229000 ;
        RECT 4.730000 0.594000 4.901000 0.649000 ;
        RECT 4.609000 0.737000 4.752000 0.792000 ;
        RECT 4.472000 0.150000 4.894000 0.205000 ;
        RECT 4.338000 0.594000 4.545000 0.649000 ;
        RECT 4.136000 0.470000 4.670000 0.525000 ;
        RECT 3.681000 0.665000 3.832000 0.720000 ;
        RECT 3.681000 0.289000 3.832000 0.344000 ;
        RECT 3.544000 0.776000 4.070000 0.831000 ;
        RECT 3.300000 0.995000 5.114000 1.050000 ;
        RECT 3.030000 0.357000 3.478000 0.412000 ;
        RECT 2.866000 0.843000 3.482000 0.898000 ;
        RECT 2.698000 0.394000 2.964000 0.449000 ;
        RECT 2.436000 0.257000 2.758000 0.312000 ;
        RECT 2.410000 0.665000 2.926000 0.720000 ;
        RECT 2.266000 0.776000 2.805000 0.831000 ;
        RECT 1.956000 0.150000 2.052000 0.205000 ;
        RECT 1.911000 0.982000 2.440000 1.037000 ;
        RECT 1.551000 0.427000 1.890000 0.482000 ;
        RECT 1.551000 0.302000 1.647000 0.357000 ;
        RECT 1.375000 0.833000 2.190000 0.888000 ;
        RECT 0.828000 0.202000 1.007000 0.257000 ;
        RECT 0.797000 0.844000 1.436000 0.899000 ;
        RECT 0.797000 0.163000 0.889000 0.218000 ;
        RECT 4.973000 0.573000 5.353000 0.627000 ;
        RECT 4.609000 0.261000 4.737000 0.315000 ;
        RECT 4.488000 0.873000 4.927000 0.927000 ;
        RECT 3.422000 0.886000 4.399000 0.940000 ;
        RECT 3.233000 0.554000 3.605000 0.608000 ;
        RECT 2.745000 0.954000 3.360000 1.008000 ;
        RECT 1.551000 0.192000 2.017000 0.246000 ;
        RECT 1.298000 0.161000 1.612000 0.215000 ;
        RECT 0.623000 0.954000 1.972000 1.008000 ;
        RECT 0.076000 0.935000 0.530000 0.989000 ;
        RECT 4.881000 0.718000 4.927000 0.927000 ;
        RECT 1.566000 0.302000 1.612000 0.749000 ;
        RECT 0.623000 0.446000 0.669000 1.008000 ;
        RECT 0.626000 0.343000 0.669000 1.008000 ;
        RECT 3.030000 0.255000 3.072000 0.650000 ;
        RECT 0.076000 0.343000 0.108000 0.989000 ;
        RECT 1.240000 0.287000 1.261000 0.738000 ;
        RECT 3.030000 0.255000 3.047000 0.783000 ;
        RECT 2.130000 0.306000 2.138000 0.902000 ;
    END
END SEDFFHQX2

MACRO SDFFSX2
    CLASS CORE ;
    FOREIGN SDFFSX2 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 4.400000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER Metal1 ;
        RECT 0.037000 0.674000 0.219000 0.767000 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.112000 0.433000 1.203000 0.595000 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 4.160000 0.694000 4.251000 0.999000 ;
        RECT 4.195000 0.177000 4.285000 0.370000 ;
        RECT 4.160000 0.694000 4.281000 0.767000 ;
        RECT 4.281000 0.315000 4.343000 0.749000 ;
        RECT 4.195000 0.315000 4.343000 0.370000 ;
        RECT 4.160000 0.694000 4.343000 0.749000 ;
        RECT 4.281000 0.177000 4.285000 0.749000 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 3.776000 0.652000 3.867000 0.733000 ;
        RECT 3.893000 0.295000 3.991000 0.361000 ;
        RECT 3.893000 0.163000 3.955000 0.707000 ;
        RECT 3.811000 0.163000 3.955000 0.218000 ;
        RECT 3.776000 0.652000 3.955000 0.707000 ;
        END
    END QN
    PIN SE
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.213000 0.433000 0.441000 0.500000 ;
        END
    END SE
    PIN SI
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.741000 0.475000 0.881000 0.633000 ;
        END
    END SI
    PIN SN
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 3.197000 0.951000 3.307000 1.033000 ;
        RECT 2.907000 0.951000 2.968000 1.026000 ;
        RECT 2.627000 0.954000 2.688000 1.026000 ;
        RECT 1.843000 0.954000 1.904000 1.010000 ;
        RECT 2.907000 0.951000 3.307000 1.006000 ;
        RECT 2.627000 0.971000 2.968000 1.026000 ;
        RECT 1.828000 0.955000 1.904000 1.010000 ;
        RECT 1.843000 0.954000 2.688000 1.008000 ;
        RECT 1.828000 0.955000 2.688000 1.008000 ;
        END
    END SN
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 4.400000 1.280000 ;
        RECT 2.384000 1.078000 2.532000 1.280000 ;
        RECT 3.968000 0.942000 4.059000 1.280000 ;
        RECT 3.440000 0.835000 3.531000 1.280000 ;
        RECT 3.045000 1.078000 3.136000 1.280000 ;
        RECT 2.048000 1.078000 2.139000 1.280000 ;
        RECT 0.853000 0.957000 0.944000 1.280000 ;
        RECT 0.197000 1.078000 0.288000 1.280000 ;
        RECT 1.675000 1.078000 1.765000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 4.400000 0.080000 ;
        RECT 2.989000 -0.080000 3.080000 0.246000 ;
        RECT 1.717000 -0.080000 1.808000 0.254000 ;
        RECT 0.865000 -0.080000 0.956000 0.122000 ;
        RECT 0.289000 -0.080000 0.380000 0.122000 ;
        RECT 3.475000 -0.080000 3.565000 0.122000 ;
        RECT 4.017000 -0.080000 4.079000 0.224000 ;
        RECT 2.340000 -0.080000 2.401000 0.328000 ;
        END
    END VSS
    OBS
        LAYER Metal1 ;
        RECT 1.268000 0.358000 1.379000 0.465000 ;
        RECT 3.248000 0.700000 3.339000 0.893000 ;
        RECT 4.037000 0.493000 4.157000 0.574000 ;
        RECT 3.653000 0.320000 3.757000 0.401000 ;
        RECT 3.632000 0.820000 3.723000 0.901000 ;
        RECT 3.492000 0.480000 3.583000 0.561000 ;
        RECT 3.331000 0.300000 3.421000 0.381000 ;
        RECT 3.312000 0.521000 3.403000 0.602000 ;
        RECT 2.908000 0.444000 2.999000 0.525000 ;
        RECT 2.723000 0.324000 2.813000 0.405000 ;
        RECT 2.485000 0.445000 2.661000 0.526000 ;
        RECT 2.251000 0.664000 2.341000 0.745000 ;
        RECT 1.632000 0.575000 1.723000 0.656000 ;
        RECT 1.441000 0.181000 1.532000 0.262000 ;
        RECT 1.391000 0.701000 1.517000 0.782000 ;
        RECT 1.228000 0.181000 1.319000 0.262000 ;
        RECT 0.940000 0.308000 1.031000 0.389000 ;
        RECT 0.568000 0.575000 0.659000 0.656000 ;
        RECT 0.544000 0.848000 0.647000 0.929000 ;
        RECT 0.503000 0.321000 0.659000 0.402000 ;
        RECT 0.411000 0.671000 0.501000 0.752000 ;
        RECT 0.048000 0.830000 0.139000 0.911000 ;
        RECT 0.048000 0.293000 0.139000 0.374000 ;
        RECT 2.095000 0.510000 2.424000 0.590000 ;
        RECT 1.917000 0.151000 2.008000 0.227000 ;
        RECT 3.653000 0.789000 3.723000 0.901000 ;
        RECT 0.048000 0.843000 0.341000 0.911000 ;
        RECT 3.312000 0.521000 3.375000 0.636000 ;
        RECT 4.037000 0.493000 4.099000 0.844000 ;
        RECT 3.653000 0.320000 3.715000 0.901000 ;
        RECT 2.937000 0.315000 2.999000 0.525000 ;
        RECT 2.485000 0.398000 2.547000 0.719000 ;
        RECT 2.217000 0.173000 2.279000 0.452000 ;
        RECT 1.661000 0.575000 1.723000 0.769000 ;
        RECT 1.005000 0.832000 1.067000 1.049000 ;
        RECT 0.597000 0.321000 0.659000 0.656000 ;
        RECT 0.585000 0.723000 0.647000 0.929000 ;
        RECT 3.492000 0.315000 3.553000 0.755000 ;
        RECT 2.751000 0.324000 2.812000 0.917000 ;
        RECT 2.623000 0.605000 2.684000 0.899000 ;
        RECT 2.095000 0.343000 2.156000 0.769000 ;
        RECT 1.787000 0.463000 1.848000 0.637000 ;
        RECT 1.604000 0.844000 1.665000 0.973000 ;
        RECT 1.456000 0.181000 1.517000 0.782000 ;
        RECT 1.399000 0.918000 1.460000 1.049000 ;
        RECT 1.268000 0.358000 1.329000 1.049000 ;
        RECT 1.132000 0.723000 1.193000 0.939000 ;
        RECT 0.731000 0.832000 0.792000 1.039000 ;
        RECT 0.643000 0.165000 0.704000 0.249000 ;
        RECT 0.440000 0.601000 0.501000 0.752000 ;
        RECT 0.388000 0.856000 0.449000 1.039000 ;
        RECT 0.280000 0.560000 0.341000 0.911000 ;
        RECT 0.048000 0.293000 0.109000 0.614000 ;
        RECT 3.653000 0.789000 4.099000 0.844000 ;
        RECT 3.248000 0.700000 3.553000 0.755000 ;
        RECT 2.937000 0.315000 3.553000 0.370000 ;
        RECT 2.751000 0.581000 3.375000 0.636000 ;
        RECT 2.251000 0.664000 2.547000 0.719000 ;
        RECT 1.787000 0.582000 2.019000 0.637000 ;
        RECT 1.661000 0.714000 2.156000 0.769000 ;
        RECT 1.604000 0.844000 2.684000 0.899000 ;
        RECT 1.532000 0.463000 1.848000 0.518000 ;
        RECT 1.517000 0.463000 1.787000 0.518000 ;
        RECT 1.456000 0.463000 1.723000 0.518000 ;
        RECT 1.399000 0.918000 1.665000 0.973000 ;
        RECT 1.005000 0.994000 1.460000 1.049000 ;
        RECT 0.731000 0.832000 1.067000 0.887000 ;
        RECT 0.643000 0.194000 1.319000 0.249000 ;
        RECT 0.503000 0.321000 1.031000 0.376000 ;
        RECT 0.503000 0.165000 0.704000 0.220000 ;
        RECT 0.440000 0.601000 0.659000 0.656000 ;
        RECT 0.048000 0.856000 0.449000 0.911000 ;
        RECT 2.217000 0.398000 2.547000 0.452000 ;
        RECT 1.917000 0.173000 2.279000 0.227000 ;
        RECT 0.585000 0.723000 1.193000 0.777000 ;
        RECT 0.388000 0.985000 0.792000 1.039000 ;
        RECT 0.048000 0.560000 0.341000 0.614000 ;
    END
END SDFFSX2

MACRO SDFFRHQX4
    CLASS CORE ;
    FOREIGN SDFFRHQX4 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 6.400000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER Metal1 ;
        RECT 0.165000 0.476000 0.290000 0.627000 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.044000 0.706000 1.206000 0.792000 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 6.091000 0.349000 6.190000 0.767000 ;
        RECT 6.244000 0.707000 6.333000 0.931000 ;
        RECT 5.918000 0.179000 6.007000 0.404000 ;
        RECT 5.573000 0.707000 5.662000 0.931000 ;
        RECT 5.540000 0.179000 5.629000 0.402000 ;
        RECT 6.244000 0.706000 6.319000 0.931000 ;
        RECT 5.555000 0.179000 5.629000 0.404000 ;
        RECT 6.091000 0.706000 6.319000 0.767000 ;
        RECT 6.091000 0.707000 6.333000 0.767000 ;
        RECT 5.573000 0.712000 6.333000 0.767000 ;
        RECT 5.555000 0.349000 6.190000 0.404000 ;
        RECT 5.540000 0.349000 6.190000 0.402000 ;
        END
    END Q
    PIN RN
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 4.529000 0.437000 4.787000 0.500000 ;
        RECT 4.527000 0.437000 4.787000 0.492000 ;
        END
    END RN
    PIN SE
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.921000 0.562000 0.981000 0.627000 ;
        RECT 0.769000 0.454000 0.829000 0.617000 ;
        RECT 0.769000 0.562000 1.090000 0.617000 ;
        RECT 0.689000 0.454000 0.829000 0.508000 ;
        END
    END SE
    PIN SI
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.729000 0.671000 0.828000 0.806000 ;
        END
    END SI
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 6.400000 1.280000 ;
        RECT 1.783000 1.078000 1.873000 1.280000 ;
        RECT 5.909000 0.910000 5.998000 1.280000 ;
        RECT 4.792000 1.078000 4.881000 1.280000 ;
        RECT 4.361000 0.989000 4.450000 1.280000 ;
        RECT 3.052000 1.078000 3.141000 1.280000 ;
        RECT 2.279000 1.078000 2.368000 1.280000 ;
        RECT 0.257000 1.078000 0.346000 1.280000 ;
        RECT 5.252000 0.742000 5.312000 1.280000 ;
        RECT 2.681000 0.982000 2.741000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 6.400000 0.080000 ;
        RECT 6.106000 -0.080000 6.196000 0.235000 ;
        RECT 1.804000 -0.080000 1.894000 0.216000 ;
        RECT 5.729000 -0.080000 5.818000 0.235000 ;
        RECT 4.834000 -0.080000 4.923000 0.122000 ;
        RECT 4.446000 -0.080000 4.535000 0.268000 ;
        RECT 2.994000 -0.080000 3.083000 0.299000 ;
        RECT 2.617000 -0.080000 2.706000 0.340000 ;
        RECT 0.962000 -0.080000 1.051000 0.122000 ;
        RECT 0.248000 -0.080000 0.337000 0.122000 ;
        RECT 5.316000 -0.080000 5.377000 0.360000 ;
        RECT 2.207000 -0.080000 2.267000 0.366000 ;
        RECT 2.192000 0.315000 2.281000 0.366000 ;
        END
    END VSS
    OBS
        LAYER Metal1 ;
        RECT 3.469000 0.285000 3.613000 0.458000 ;
        RECT 2.053000 0.699000 2.443000 0.792000 ;
        RECT 1.900000 0.480000 1.993000 0.615000 ;
        RECT 0.043000 0.729000 0.136000 0.952000 ;
        RECT 0.043000 0.167000 0.136000 0.360000 ;
        RECT 3.712000 0.161000 3.801000 0.329000 ;
        RECT 5.196000 0.506000 5.314000 0.594000 ;
        RECT 2.018000 0.294000 2.116000 0.381000 ;
        RECT 1.001000 0.344000 1.090000 0.431000 ;
        RECT 1.512000 0.480000 1.616000 0.563000 ;
        RECT 4.635000 0.236000 4.724000 0.317000 ;
        RECT 4.083000 0.262000 4.179000 0.343000 ;
        RECT 2.806000 0.270000 2.895000 0.351000 ;
        RECT 2.650000 0.655000 2.739000 0.736000 ;
        RECT 1.924000 0.698000 2.116000 0.779000 ;
        RECT 1.726000 0.612000 1.815000 0.693000 ;
        RECT 1.549000 0.650000 1.638000 0.731000 ;
        RECT 1.498000 0.214000 1.587000 0.295000 ;
        RECT 0.455000 0.476000 0.544000 0.557000 ;
        RECT 0.605000 0.208000 0.695000 0.287000 ;
        RECT 4.010000 0.627000 4.143000 0.704000 ;
        RECT 4.649000 0.192000 4.724000 0.317000 ;
        RECT 3.474000 0.692000 3.549000 0.792000 ;
        RECT 1.309000 0.208000 1.401000 0.275000 ;
        RECT 2.053000 0.698000 2.116000 0.792000 ;
        RECT 4.231000 0.862000 4.292000 1.039000 ;
        RECT 3.488000 0.285000 3.549000 0.792000 ;
        RECT 3.353000 0.815000 3.414000 0.915000 ;
        RECT 3.336000 0.421000 3.397000 0.580000 ;
        RECT 3.201000 0.954000 3.262000 1.039000 ;
        RECT 3.197000 0.285000 3.258000 0.425000 ;
        RECT 2.834000 0.270000 2.895000 0.425000 ;
        RECT 2.247000 0.919000 2.308000 0.994000 ;
        RECT 1.563000 0.650000 1.624000 0.994000 ;
        RECT 1.424000 0.508000 1.485000 0.818000 ;
        RECT 1.386000 0.350000 1.447000 0.437000 ;
        RECT 0.043000 0.167000 0.104000 0.952000 ;
        RECT 5.196000 0.192000 5.256000 0.594000 ;
        RECT 5.132000 0.539000 5.192000 0.994000 ;
        RECT 5.075000 0.301000 5.135000 0.423000 ;
        RECT 5.011000 0.524000 5.071000 0.885000 ;
        RECT 4.884000 0.368000 4.944000 0.775000 ;
        RECT 4.647000 0.751000 4.707000 0.885000 ;
        RECT 4.513000 0.862000 4.573000 0.994000 ;
        RECT 4.407000 0.524000 4.467000 0.665000 ;
        RECT 4.285000 0.649000 4.345000 0.806000 ;
        RECT 4.111000 0.762000 4.171000 0.915000 ;
        RECT 4.083000 0.161000 4.143000 0.704000 ;
        RECT 3.863000 0.285000 3.923000 0.458000 ;
        RECT 3.626000 0.600000 3.686000 0.682000 ;
        RECT 3.057000 0.660000 3.117000 0.746000 ;
        RECT 2.922000 0.525000 2.982000 0.870000 ;
        RECT 2.802000 0.808000 2.862000 1.008000 ;
        RECT 2.664000 0.423000 2.724000 0.736000 ;
        RECT 2.542000 0.919000 2.602000 1.005000 ;
        RECT 2.504000 0.546000 2.564000 0.863000 ;
        RECT 2.456000 0.300000 2.516000 0.477000 ;
        RECT 2.427000 0.161000 2.487000 0.381000 ;
        RECT 2.056000 0.294000 2.116000 0.792000 ;
        RECT 1.755000 0.612000 1.815000 0.752000 ;
        RECT 1.512000 0.214000 1.572000 0.563000 ;
        RECT 1.266000 0.382000 1.326000 0.932000 ;
        RECT 0.607000 0.775000 0.667000 0.932000 ;
        RECT 0.485000 0.885000 0.545000 1.042000 ;
        RECT 0.469000 0.256000 0.529000 0.720000 ;
        RECT 1.266000 0.874000 1.624000 0.932000 ;
        RECT 5.196000 0.506000 5.902000 0.561000 ;
        RECT 5.132000 0.539000 5.314000 0.594000 ;
        RECT 4.884000 0.368000 5.135000 0.423000 ;
        RECT 4.647000 0.830000 5.071000 0.885000 ;
        RECT 4.513000 0.939000 5.192000 0.994000 ;
        RECT 4.285000 0.751000 4.707000 0.806000 ;
        RECT 4.252000 0.524000 4.467000 0.579000 ;
        RECT 4.231000 0.862000 4.573000 0.917000 ;
        RECT 4.010000 0.649000 4.345000 0.704000 ;
        RECT 3.626000 0.627000 4.143000 0.682000 ;
        RECT 3.474000 0.737000 3.900000 0.792000 ;
        RECT 2.922000 0.815000 3.414000 0.870000 ;
        RECT 2.834000 0.370000 3.258000 0.425000 ;
        RECT 2.664000 0.525000 3.397000 0.580000 ;
        RECT 2.504000 0.808000 2.862000 0.863000 ;
        RECT 2.247000 0.919000 2.602000 0.974000 ;
        RECT 2.177000 0.546000 2.564000 0.601000 ;
        RECT 1.563000 0.939000 2.308000 0.994000 ;
        RECT 1.512000 0.480000 1.993000 0.535000 ;
        RECT 1.424000 0.508000 1.616000 0.563000 ;
        RECT 1.266000 0.382000 1.447000 0.437000 ;
        RECT 0.607000 0.877000 1.624000 0.932000 ;
        RECT 0.605000 0.208000 1.401000 0.263000 ;
        RECT 0.485000 0.987000 1.300000 1.042000 ;
        RECT 0.469000 0.344000 1.090000 0.399000 ;
        RECT 0.440000 0.665000 0.529000 0.720000 ;
        RECT 0.422000 0.256000 0.529000 0.311000 ;
        RECT 0.043000 0.775000 0.667000 0.830000 ;
        RECT 4.649000 0.192000 5.256000 0.246000 ;
        RECT 4.407000 0.611000 4.944000 0.665000 ;
        RECT 3.863000 0.285000 3.990000 0.339000 ;
        RECT 3.469000 0.404000 3.923000 0.458000 ;
        RECT 3.353000 0.861000 4.171000 0.915000 ;
        RECT 3.324000 0.161000 4.143000 0.215000 ;
        RECT 3.201000 0.985000 4.292000 1.039000 ;
        RECT 3.197000 0.285000 3.613000 0.339000 ;
        RECT 3.057000 0.692000 3.549000 0.746000 ;
        RECT 2.802000 0.954000 3.262000 1.008000 ;
        RECT 2.456000 0.423000 2.724000 0.477000 ;
        RECT 2.331000 0.161000 2.487000 0.215000 ;
        RECT 1.755000 0.698000 2.116000 0.752000 ;
        RECT 0.451000 0.885000 0.545000 0.939000 ;
        RECT 2.456000 0.161000 2.487000 0.477000 ;
    END
END SDFFRHQX4

MACRO SDFFRHQX2
    CLASS CORE ;
    FOREIGN SDFFRHQX2 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 5.200000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER Metal1 ;
        RECT 0.158000 0.506000 0.310000 0.617000 ;
        RECT 0.230000 0.506000 0.290000 0.627000 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.019000 0.418000 1.177000 0.510000 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 4.551000 0.225000 4.643000 0.330000 ;
        RECT 4.727000 0.674000 4.817000 0.960000 ;
        RECT 4.551000 0.151000 4.641000 0.344000 ;
        RECT 4.937000 0.275000 4.998000 0.729000 ;
        RECT 4.727000 0.674000 4.998000 0.729000 ;
        RECT 4.551000 0.275000 4.998000 0.330000 ;
        END
    END Q
    PIN RN
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 4.216000 0.632000 4.357000 0.763000 ;
        END
    END RN
    PIN SE
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.383000 0.415000 0.491000 0.543000 ;
        END
    END SE
    PIN SI
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.776000 0.548000 0.865000 0.629000 ;
        RECT 0.776000 0.567000 0.984000 0.629000 ;
        END
    END SI
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 5.200000 1.280000 ;
        RECT 3.662000 1.078000 3.778000 1.280000 ;
        RECT 0.236000 1.013000 0.347000 1.280000 ;
        RECT 5.063000 0.800000 5.153000 1.280000 ;
        RECT 4.367000 1.078000 4.457000 1.280000 ;
        RECT 4.000000 1.078000 4.089000 1.280000 ;
        RECT 2.670000 1.078000 2.759000 1.280000 ;
        RECT 1.665000 0.997000 1.754000 1.280000 ;
        RECT 0.830000 1.001000 0.919000 1.280000 ;
        RECT 0.247000 0.972000 0.336000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 4.135000 -0.080000 4.382000 0.122000 ;
        RECT 0.000000 -0.080000 5.200000 0.080000 ;
        RECT 2.664000 -0.080000 2.754000 0.292000 ;
        RECT 1.641000 -0.080000 1.731000 0.327000 ;
        RECT 0.194000 -0.080000 0.284000 0.122000 ;
        RECT 4.751000 -0.080000 4.840000 0.122000 ;
        RECT 3.693000 -0.080000 3.782000 0.122000 ;
        RECT 0.737000 -0.080000 0.826000 0.122000 ;
        RECT 1.670000 -0.080000 1.731000 0.328000 ;
        END
    END VSS
    OBS
        LAYER Metal1 ;
        RECT 3.058000 0.206000 3.158000 0.419000 ;
        RECT 1.359000 0.698000 1.454000 0.792000 ;
        RECT 3.334000 0.170000 3.425000 0.261000 ;
        RECT 4.199000 0.352000 4.289000 0.577000 ;
        RECT 2.853000 0.240000 2.943000 0.417000 ;
        RECT 1.825000 0.398000 1.915000 0.532000 ;
        RECT 0.047000 0.671000 0.137000 0.864000 ;
        RECT 4.473000 0.523000 4.562000 0.612000 ;
        RECT 1.743000 0.607000 1.832000 0.701000 ;
        RECT 0.552000 0.323000 0.852000 0.405000 ;
        RECT 4.664000 0.538000 4.877000 0.619000 ;
        RECT 4.226000 0.838000 4.315000 0.919000 ;
        RECT 4.005000 0.517000 4.094000 0.598000 ;
        RECT 3.921000 0.336000 4.010000 0.417000 ;
        RECT 3.732000 0.736000 3.821000 0.817000 ;
        RECT 3.658000 0.605000 3.807000 0.686000 ;
        RECT 3.369000 0.633000 3.459000 0.714000 ;
        RECT 3.245000 0.795000 3.362000 0.876000 ;
        RECT 3.236000 0.338000 3.325000 0.419000 ;
        RECT 2.894000 0.804000 2.983000 0.885000 ;
        RECT 2.532000 0.802000 2.621000 0.883000 ;
        RECT 2.348000 0.748000 2.437000 0.829000 ;
        RECT 2.247000 0.293000 2.336000 0.374000 ;
        RECT 1.853000 0.795000 1.976000 0.876000 ;
        RECT 1.812000 0.150000 1.901000 0.231000 ;
        RECT 1.419000 0.902000 1.509000 0.983000 ;
        RECT 1.283000 0.150000 1.372000 0.231000 ;
        RECT 1.098000 0.202000 1.187000 0.283000 ;
        RECT 0.599000 0.595000 0.688000 0.676000 ;
        RECT 0.552000 0.324000 0.901000 0.405000 ;
        RECT 0.525000 0.938000 0.615000 1.019000 ;
        RECT 0.047000 0.318000 0.137000 0.399000 ;
        RECT 3.409000 0.360000 3.498000 0.440000 ;
        RECT 1.567000 0.510000 1.656000 0.590000 ;
        RECT 3.732000 0.605000 3.807000 0.817000 ;
        RECT 1.419000 0.901000 1.494000 0.983000 ;
        RECT 0.047000 0.318000 0.122000 0.450000 ;
        RECT 0.552000 0.323000 0.624000 0.663000 ;
        RECT 3.832000 0.206000 3.925000 0.273000 ;
        RECT 3.245000 0.795000 3.310000 0.915000 ;
        RECT 4.664000 0.399000 4.725000 0.619000 ;
        RECT 4.350000 0.206000 4.411000 0.454000 ;
        RECT 3.964000 0.543000 4.025000 0.994000 ;
        RECT 3.746000 0.349000 3.807000 0.817000 ;
        RECT 3.423000 0.360000 3.484000 0.688000 ;
        RECT 2.907000 0.362000 2.968000 0.885000 ;
        RECT 2.786000 0.471000 2.847000 0.746000 ;
        RECT 2.123000 0.607000 2.184000 0.994000 ;
        RECT 1.595000 0.477000 1.656000 0.590000 ;
        RECT 1.393000 0.176000 1.454000 0.792000 ;
        RECT 1.238000 0.575000 1.299000 0.956000 ;
        RECT 1.117000 0.856000 1.178000 0.995000 ;
        RECT 0.538000 0.732000 0.599000 0.858000 ;
        RECT 0.408000 0.608000 0.469000 0.748000 ;
        RECT 3.371000 0.939000 3.431000 1.039000 ;
        RECT 3.245000 0.338000 3.305000 0.915000 ;
        RECT 3.098000 0.206000 3.158000 0.786000 ;
        RECT 2.977000 0.817000 3.037000 0.915000 ;
        RECT 2.856000 0.939000 2.916000 1.039000 ;
        RECT 2.490000 0.252000 2.550000 0.417000 ;
        RECT 2.377000 0.692000 2.437000 0.829000 ;
        RECT 2.368000 0.319000 2.428000 0.526000 ;
        RECT 2.247000 0.477000 2.307000 0.637000 ;
        RECT 2.247000 0.176000 2.307000 0.374000 ;
        RECT 1.916000 0.477000 1.976000 0.876000 ;
        RECT 1.241000 0.445000 1.301000 0.630000 ;
        RECT 0.695000 0.856000 0.755000 0.993000 ;
        RECT 0.485000 0.165000 0.545000 0.261000 ;
        RECT 0.037000 0.395000 0.097000 0.726000 ;
        RECT 1.241000 0.445000 1.299000 0.956000 ;
        RECT 4.350000 0.399000 4.725000 0.454000 ;
        RECT 3.964000 0.838000 4.315000 0.893000 ;
        RECT 3.746000 0.349000 4.010000 0.404000 ;
        RECT 3.371000 0.939000 4.025000 0.994000 ;
        RECT 3.058000 0.206000 4.411000 0.261000 ;
        RECT 2.490000 0.362000 2.968000 0.417000 ;
        RECT 2.368000 0.471000 2.847000 0.526000 ;
        RECT 2.247000 0.582000 2.684000 0.637000 ;
        RECT 2.247000 0.319000 2.428000 0.374000 ;
        RECT 2.123000 0.939000 2.916000 0.994000 ;
        RECT 1.812000 0.176000 2.307000 0.231000 ;
        RECT 1.595000 0.477000 2.307000 0.532000 ;
        RECT 1.393000 0.646000 1.832000 0.701000 ;
        RECT 1.283000 0.176000 1.454000 0.231000 ;
        RECT 1.238000 0.901000 1.494000 0.956000 ;
        RECT 0.695000 0.856000 1.178000 0.911000 ;
        RECT 0.538000 0.732000 1.299000 0.787000 ;
        RECT 0.525000 0.938000 0.755000 0.993000 ;
        RECT 0.485000 0.206000 1.187000 0.261000 ;
        RECT 0.408000 0.608000 0.688000 0.663000 ;
        RECT 0.378000 0.165000 0.545000 0.220000 ;
        RECT 4.005000 0.523000 4.562000 0.577000 ;
        RECT 2.977000 0.861000 3.310000 0.915000 ;
        RECT 2.856000 0.985000 3.431000 1.039000 ;
        RECT 2.532000 0.817000 3.037000 0.871000 ;
        RECT 2.377000 0.692000 2.847000 0.746000 ;
        RECT 0.047000 0.804000 0.599000 0.858000 ;
        RECT 0.047000 0.318000 0.097000 0.864000 ;
        RECT 3.423000 0.360000 3.459000 0.714000 ;
        RECT 2.907000 0.240000 2.943000 0.885000 ;
        RECT 0.599000 0.323000 0.624000 0.676000 ;
        RECT 4.005000 0.517000 4.025000 0.994000 ;
        RECT 2.977000 0.804000 2.983000 0.915000 ;
    END
END SDFFRHQX2

MACRO SDFFRX2
    CLASS CORE ;
    FOREIGN SDFFRX2 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 5.200000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER Metal1 ;
        RECT 0.164000 0.408000 0.253000 0.671000 ;
        RECT 0.164000 0.429000 0.302000 0.505000 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.008000 0.369000 1.177000 0.505000 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 5.050000 0.227000 5.159000 0.387000 ;
        RECT 5.050000 0.163000 5.140000 0.387000 ;
        RECT 5.053000 0.693000 5.142000 0.779000 ;
        RECT 5.045000 0.698000 5.142000 0.779000 ;
        RECT 5.081000 0.227000 5.159000 0.769000 ;
        RECT 5.053000 0.693000 5.159000 0.769000 ;
        RECT 5.045000 0.698000 5.159000 0.769000 ;
        RECT 5.081000 0.227000 5.142000 0.779000 ;
        RECT 5.081000 0.163000 5.140000 0.779000 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 4.706000 0.698000 4.796000 0.779000 ;
        RECT 4.643000 0.326000 4.733000 0.407000 ;
        RECT 4.672000 0.326000 4.733000 0.489000 ;
        RECT 4.721000 0.435000 4.781000 0.779000 ;
        RECT 4.721000 0.435000 4.797000 0.494000 ;
        RECT 4.672000 0.435000 4.797000 0.489000 ;
        RECT 4.721000 0.326000 4.733000 0.779000 ;
        END
    END QN
    PIN RN
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.790000 0.656000 1.903000 0.794000 ;
        RECT 1.790000 0.685000 1.917000 0.794000 ;
        RECT 1.828000 0.685000 1.917000 0.807000 ;
        RECT 1.778000 0.685000 1.917000 0.771000 ;
        RECT 1.828000 0.656000 1.903000 0.807000 ;
        END
    END RN
    PIN SE
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.376000 0.460000 0.465000 0.540000 ;
        RECT 0.390000 0.295000 0.471000 0.371000 ;
        RECT 0.390000 0.295000 0.450000 0.540000 ;
        END
    END SE
    PIN SI
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.743000 0.538000 0.902000 0.638000 ;
        END
    END SI
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 2.600000 1.047000 2.979000 1.280000 ;
        RECT 0.000000 1.120000 5.200000 1.280000 ;
        RECT 4.874000 0.986000 4.964000 1.280000 ;
        RECT 4.333000 0.891000 4.423000 1.280000 ;
        RECT 3.603000 0.986000 3.693000 1.280000 ;
        RECT 0.194000 1.078000 0.284000 1.280000 ;
        RECT 1.749000 1.078000 1.838000 1.280000 ;
        RECT 0.919000 0.963000 1.008000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 1.926000 -0.080000 2.358000 0.090000 ;
        RECT 0.000000 -0.080000 5.200000 0.080000 ;
        RECT 1.926000 -0.080000 2.038000 0.303000 ;
        RECT 4.312000 -0.080000 4.402000 0.268000 ;
        RECT 0.735000 -0.080000 0.825000 0.122000 ;
        RECT 0.194000 -0.080000 0.284000 0.122000 ;
        RECT 3.921000 -0.080000 4.010000 0.122000 ;
        RECT 3.433000 -0.080000 3.522000 0.283000 ;
        RECT 2.716000 -0.080000 2.805000 0.311000 ;
        RECT 2.269000 -0.080000 2.358000 0.214000 ;
        RECT 4.860000 -0.080000 4.920000 0.355000 ;
        END
    END VSS
    OBS
        LAYER Metal1 ;
        RECT 3.616000 0.292000 3.737000 0.418000 ;
        RECT 3.761000 0.638000 3.858000 0.794000 ;
        RECT 3.763000 0.586000 3.858000 0.794000 ;
        RECT 1.891000 0.483000 2.035000 0.577000 ;
        RECT 0.043000 0.864000 0.137000 1.008000 ;
        RECT 4.522000 0.851000 4.612000 0.957000 ;
        RECT 4.373000 0.379000 4.462000 0.487000 ;
        RECT 2.847000 0.517000 2.936000 0.687000 ;
        RECT 1.765000 0.161000 1.854000 0.264000 ;
        RECT 1.093000 0.206000 1.182000 0.302000 ;
        RECT 0.544000 0.348000 0.633000 0.493000 ;
        RECT 1.573000 0.373000 1.660000 0.496000 ;
        RECT 4.512000 0.158000 4.601000 0.239000 ;
        RECT 4.123000 0.217000 4.213000 0.298000 ;
        RECT 3.950000 0.781000 4.039000 0.862000 ;
        RECT 3.884000 0.388000 3.974000 0.469000 ;
        RECT 3.876000 0.936000 4.010000 1.017000 ;
        RECT 3.763000 0.586000 3.989000 0.667000 ;
        RECT 3.257000 0.774000 3.346000 0.855000 ;
        RECT 3.194000 0.619000 3.283000 0.700000 ;
        RECT 2.671000 0.626000 2.760000 0.707000 ;
        RECT 2.235000 0.826000 2.324000 0.907000 ;
        RECT 2.138000 0.346000 2.227000 0.427000 ;
        RECT 2.022000 0.845000 2.112000 0.926000 ;
        RECT 1.571000 0.415000 1.660000 0.496000 ;
        RECT 1.418000 0.786000 1.507000 0.867000 ;
        RECT 1.303000 0.221000 1.488000 0.302000 ;
        RECT 1.276000 0.945000 1.366000 1.026000 ;
        RECT 1.238000 0.381000 1.328000 0.462000 ;
        RECT 1.104000 0.679000 1.194000 0.760000 ;
        RECT 0.793000 0.389000 0.882000 0.470000 ;
        RECT 0.404000 0.817000 0.494000 0.898000 ;
        RECT 0.043000 0.262000 0.137000 0.343000 ;
        RECT 3.073000 0.260000 3.178000 0.340000 ;
        RECT 2.210000 0.510000 2.299000 0.590000 ;
        RECT 2.519000 0.287000 2.595000 0.461000 ;
        RECT 3.899000 0.388000 3.974000 0.487000 ;
        RECT 2.519000 0.274000 2.593000 0.461000 ;
        RECT 0.378000 0.158000 0.469000 0.229000 ;
        RECT 2.570000 0.639000 2.760000 0.707000 ;
        RECT 1.427000 0.781000 1.493000 0.867000 ;
        RECT 4.887000 0.577000 4.948000 0.906000 ;
        RECT 4.522000 0.158000 4.583000 0.957000 ;
        RECT 4.387000 0.379000 4.448000 0.754000 ;
        RECT 4.152000 0.217000 4.213000 0.487000 ;
        RECT 3.763000 0.401000 3.824000 0.794000 ;
        RECT 3.465000 0.473000 3.526000 0.581000 ;
        RECT 3.129000 0.645000 3.190000 0.929000 ;
        RECT 3.117000 0.260000 3.178000 0.418000 ;
        RECT 2.504000 0.158000 2.565000 0.355000 ;
        RECT 2.454000 0.874000 2.515000 1.037000 ;
        RECT 2.249000 0.704000 2.310000 0.907000 ;
        RECT 1.900000 0.939000 1.961000 1.037000 ;
        RECT 1.427000 0.161000 1.488000 0.867000 ;
        RECT 1.091000 0.821000 1.152000 1.000000 ;
        RECT 0.613000 0.158000 0.674000 0.261000 ;
        RECT 0.600000 0.821000 0.661000 1.008000 ;
        RECT 0.525000 0.438000 0.586000 0.652000 ;
        RECT 0.433000 0.676000 0.494000 0.898000 ;
        RECT 0.043000 0.262000 0.104000 1.008000 ;
        RECT 4.960000 0.455000 5.020000 0.632000 ;
        RECT 4.184000 0.699000 4.244000 0.836000 ;
        RECT 3.950000 0.781000 4.010000 1.017000 ;
        RECT 3.677000 0.292000 3.737000 0.456000 ;
        RECT 3.434000 0.739000 3.494000 0.829000 ;
        RECT 2.997000 0.406000 3.057000 0.818000 ;
        RECT 2.570000 0.639000 2.630000 0.929000 ;
        RECT 2.360000 0.375000 2.420000 0.758000 ;
        RECT 2.167000 0.346000 2.227000 0.430000 ;
        RECT 2.037000 0.523000 2.097000 0.926000 ;
        RECT 1.606000 0.939000 1.666000 1.013000 ;
        RECT 1.279000 0.394000 1.339000 1.026000 ;
        RECT 0.482000 0.596000 0.542000 0.757000 ;
        RECT 3.628000 0.525000 3.689000 0.581000 ;
        RECT 4.887000 0.577000 5.020000 0.632000 ;
        RECT 4.522000 0.851000 4.948000 0.906000 ;
        RECT 4.184000 0.699000 4.448000 0.754000 ;
        RECT 3.950000 0.781000 4.244000 0.836000 ;
        RECT 3.899000 0.432000 4.462000 0.487000 ;
        RECT 3.677000 0.401000 3.824000 0.456000 ;
        RECT 3.628000 0.525000 3.703000 0.580000 ;
        RECT 3.465000 0.526000 3.689000 0.581000 ;
        RECT 3.434000 0.739000 3.858000 0.794000 ;
        RECT 3.257000 0.774000 3.494000 0.829000 ;
        RECT 3.129000 0.645000 3.283000 0.700000 ;
        RECT 3.117000 0.363000 3.737000 0.418000 ;
        RECT 2.750000 0.763000 3.057000 0.818000 ;
        RECT 2.519000 0.406000 3.057000 0.461000 ;
        RECT 2.454000 0.874000 3.190000 0.929000 ;
        RECT 2.435000 0.158000 2.565000 0.213000 ;
        RECT 2.167000 0.375000 2.420000 0.430000 ;
        RECT 1.900000 0.982000 2.515000 1.037000 ;
        RECT 1.606000 0.939000 1.961000 0.994000 ;
        RECT 1.276000 0.958000 1.666000 1.013000 ;
        RECT 1.091000 0.945000 1.366000 1.000000 ;
        RECT 0.650000 0.699000 1.194000 0.754000 ;
        RECT 0.613000 0.206000 1.182000 0.261000 ;
        RECT 0.600000 0.821000 1.152000 0.876000 ;
        RECT 0.544000 0.402000 0.882000 0.457000 ;
        RECT 0.378000 0.158000 0.674000 0.213000 ;
        RECT 2.997000 0.473000 3.526000 0.527000 ;
        RECT 2.360000 0.517000 2.936000 0.571000 ;
        RECT 2.249000 0.704000 2.420000 0.758000 ;
        RECT 1.891000 0.523000 2.299000 0.577000 ;
        RECT 1.573000 0.373000 2.227000 0.427000 ;
        RECT 1.427000 0.161000 1.854000 0.215000 ;
        RECT 0.043000 0.954000 0.661000 1.008000 ;
        RECT 1.279000 0.381000 1.328000 1.026000 ;
        RECT 2.519000 0.158000 2.565000 0.461000 ;
        RECT 0.544000 0.348000 0.586000 0.652000 ;
        RECT 0.525000 0.438000 0.542000 0.757000 ;
        RECT 0.482000 0.596000 0.494000 0.898000 ;
    END
END SDFFRX2

MACRO SDFFHQX4
    CLASS CORE ;
    FOREIGN SDFFHQX4 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 4.500000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER Metal1 ;
        RECT 0.152000 0.524000 0.290000 0.627000 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.067000 0.356000 1.156000 0.437000 ;
        RECT 1.088000 0.356000 1.156000 0.439000 ;
        RECT 1.088000 0.356000 1.150000 0.627000 ;
        RECT 1.088000 0.573000 1.155000 0.627000 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 4.191000 0.433000 4.290000 0.767000 ;
        RECT 4.193000 0.325000 4.282000 0.767000 ;
        RECT 4.130000 0.671000 4.290000 0.752000 ;
        END
    END Q
    PIN SE
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.926000 0.593000 1.015000 0.674000 ;
        RECT 0.527000 0.567000 0.690000 0.633000 ;
        RECT 0.629000 0.567000 0.690000 0.656000 ;
        RECT 0.629000 0.601000 1.015000 0.656000 ;
        END
    END SE
    PIN SI
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.750000 0.433000 0.871000 0.533000 ;
        RECT 0.750000 0.433000 0.839000 0.546000 ;
        RECT 0.729000 0.433000 0.871000 0.500000 ;
        END
    END SI
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 3.060000 1.078000 3.687000 1.280000 ;
        RECT 0.000000 1.120000 4.500000 1.280000 ;
        RECT 4.299000 0.989000 4.389000 1.280000 ;
        RECT 3.951000 1.078000 4.040000 1.280000 ;
        RECT 2.284000 1.078000 2.373000 1.280000 ;
        RECT 1.390000 1.078000 1.479000 1.280000 ;
        RECT 0.248000 1.078000 0.337000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 4.500000 0.080000 ;
        RECT 4.025000 -0.080000 4.115000 0.212000 ;
        RECT 4.361000 -0.080000 4.450000 0.215000 ;
        RECT 3.632000 -0.080000 3.721000 0.122000 ;
        RECT 1.678000 -0.080000 1.767000 0.287000 ;
        RECT 0.755000 -0.080000 0.844000 0.122000 ;
        RECT 0.249000 -0.080000 0.338000 0.410000 ;
        RECT 2.361000 -0.080000 2.422000 0.311000 ;
        RECT 3.185000 -0.080000 3.245000 0.287000 ;
        RECT 0.249000 0.359000 0.346000 0.410000 ;
        END
    END VSS
    OBS
        LAYER Metal1 ;
        RECT 0.399000 0.154000 0.490000 0.246000 ;
        RECT 0.490000 0.318000 0.580000 0.425000 ;
        RECT 3.380000 0.150000 3.469000 0.412000 ;
        RECT 2.596000 0.605000 2.685000 0.787000 ;
        RECT 0.047000 0.739000 0.136000 0.932000 ;
        RECT 0.406000 0.692000 0.509000 0.779000 ;
        RECT 1.112000 0.160000 1.201000 0.246000 ;
        RECT 3.842000 0.264000 3.931000 0.345000 ;
        RECT 3.842000 0.264000 3.923000 0.571000 ;
        RECT 3.799000 0.826000 3.923000 0.907000 ;
        RECT 3.699000 0.490000 3.923000 0.571000 ;
        RECT 3.576000 0.650000 3.802000 0.731000 ;
        RECT 3.265000 0.577000 3.354000 0.658000 ;
        RECT 2.913000 0.348000 3.003000 0.429000 ;
        RECT 2.911000 0.596000 3.000000 0.677000 ;
        RECT 2.725000 0.223000 2.814000 0.304000 ;
        RECT 2.672000 0.954000 2.761000 1.035000 ;
        RECT 2.536000 0.245000 2.628000 0.326000 ;
        RECT 2.483000 0.843000 2.573000 0.924000 ;
        RECT 2.420000 0.490000 2.510000 0.571000 ;
        RECT 2.221000 0.504000 2.310000 0.585000 ;
        RECT 2.137000 0.789000 2.226000 0.870000 ;
        RECT 2.010000 0.454000 2.161000 0.535000 ;
        RECT 1.952000 0.790000 2.042000 0.871000 ;
        RECT 1.867000 0.273000 1.956000 0.354000 ;
        RECT 1.740000 0.450000 1.829000 0.531000 ;
        RECT 1.689000 0.612000 1.950000 0.693000 ;
        RECT 1.545000 0.938000 1.634000 1.019000 ;
        RECT 1.248000 0.331000 1.337000 0.412000 ;
        RECT 1.193000 0.776000 1.282000 0.857000 ;
        RECT 0.606000 0.724000 0.695000 0.805000 ;
        RECT 0.068000 0.344000 0.157000 0.425000 ;
        RECT 0.047000 0.688000 0.122000 0.932000 ;
        RECT 1.889000 0.790000 2.042000 0.858000 ;
        RECT 3.414000 0.467000 3.475000 0.768000 ;
        RECT 3.064000 0.223000 3.125000 0.412000 ;
        RECT 3.060000 0.604000 3.121000 0.787000 ;
        RECT 2.942000 0.348000 3.003000 0.521000 ;
        RECT 2.567000 0.245000 2.628000 0.429000 ;
        RECT 2.420000 0.381000 2.481000 0.571000 ;
        RECT 2.137000 0.679000 2.198000 0.870000 ;
        RECT 2.120000 0.269000 2.181000 0.402000 ;
        RECT 1.889000 0.273000 1.950000 0.858000 ;
        RECT 1.463000 0.163000 1.524000 0.855000 ;
        RECT 1.084000 0.939000 1.145000 1.050000 ;
        RECT 0.490000 0.318000 0.551000 0.512000 ;
        RECT 0.422000 0.877000 0.483000 1.050000 ;
        RECT 0.406000 0.457000 0.467000 0.779000 ;
        RECT 0.031000 0.369000 0.092000 0.743000 ;
        RECT 3.863000 0.264000 3.923000 0.907000 ;
        RECT 3.576000 0.357000 3.636000 0.886000 ;
        RECT 3.303000 0.831000 3.363000 1.008000 ;
        RECT 3.181000 0.713000 3.241000 0.898000 ;
        RECT 2.747000 0.490000 2.807000 0.652000 ;
        RECT 2.287000 0.530000 2.347000 0.993000 ;
        RECT 2.241000 0.158000 2.301000 0.436000 ;
        RECT 2.101000 0.348000 2.161000 0.733000 ;
        RECT 1.896000 0.158000 1.956000 0.354000 ;
        RECT 1.343000 0.357000 1.403000 0.994000 ;
        RECT 0.952000 0.802000 1.012000 0.936000 ;
        RECT 0.031000 0.369000 0.157000 0.425000 ;
        RECT 3.303000 0.831000 3.636000 0.886000 ;
        RECT 3.181000 0.713000 3.475000 0.768000 ;
        RECT 3.064000 0.357000 3.636000 0.412000 ;
        RECT 2.567000 0.374000 3.003000 0.429000 ;
        RECT 2.483000 0.843000 3.241000 0.898000 ;
        RECT 2.483000 0.490000 2.807000 0.545000 ;
        RECT 2.420000 0.490000 2.725000 0.545000 ;
        RECT 2.287000 0.732000 3.121000 0.787000 ;
        RECT 2.241000 0.381000 2.481000 0.436000 ;
        RECT 2.221000 0.530000 2.347000 0.585000 ;
        RECT 1.896000 0.158000 2.301000 0.213000 ;
        RECT 1.545000 0.938000 2.347000 0.993000 ;
        RECT 1.545000 0.450000 1.829000 0.505000 ;
        RECT 1.524000 0.450000 1.740000 0.505000 ;
        RECT 1.463000 0.450000 1.689000 0.505000 ;
        RECT 1.322000 0.163000 1.524000 0.218000 ;
        RECT 1.248000 0.357000 1.403000 0.412000 ;
        RECT 1.084000 0.939000 1.634000 0.994000 ;
        RECT 0.952000 0.802000 1.282000 0.857000 ;
        RECT 0.543000 0.881000 1.012000 0.936000 ;
        RECT 0.490000 0.318000 0.952000 0.373000 ;
        RECT 0.422000 0.995000 1.145000 1.050000 ;
        RECT 0.406000 0.724000 0.695000 0.779000 ;
        RECT 0.406000 0.457000 0.551000 0.512000 ;
        RECT 0.047000 0.877000 0.483000 0.932000 ;
        RECT 0.031000 0.688000 0.122000 0.743000 ;
        RECT 3.060000 0.604000 3.354000 0.658000 ;
        RECT 2.942000 0.467000 3.475000 0.521000 ;
        RECT 2.747000 0.598000 3.000000 0.652000 ;
        RECT 2.725000 0.223000 3.125000 0.277000 ;
        RECT 2.672000 0.954000 3.363000 1.008000 ;
        RECT 2.101000 0.679000 2.198000 0.733000 ;
        RECT 2.101000 0.348000 2.181000 0.402000 ;
        RECT 1.896000 0.158000 1.950000 0.858000 ;
        RECT 1.084000 0.939000 2.347000 0.993000 ;
        RECT 0.399000 0.192000 1.201000 0.246000 ;
        RECT 2.137000 0.269000 2.161000 0.870000 ;
        RECT 0.068000 0.344000 0.092000 0.932000 ;
        RECT 2.287000 0.504000 2.310000 0.993000 ;
        RECT 0.047000 0.369000 0.068000 0.932000 ;
        RECT 2.120000 0.269000 2.137000 0.733000 ;
    END
END SDFFHQX4

MACRO SDFFHQX2
    CLASS CORE ;
    FOREIGN SDFFHQX2 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 4.200000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER Metal1 ;
        RECT 0.212000 0.512000 0.327000 0.633000 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.051000 0.335000 1.184000 0.494000 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 3.855000 0.167000 3.945000 0.248000 ;
        RECT 3.695000 0.700000 3.813000 0.767000 ;
        RECT 3.695000 0.193000 3.756000 0.767000 ;
        RECT 3.695000 0.193000 3.945000 0.248000 ;
        END
    END Q
    PIN SE
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.998000 0.648000 1.088000 0.729000 ;
        RECT 0.562000 0.567000 0.663000 0.635000 ;
        RECT 0.544000 0.568000 0.663000 0.635000 ;
        RECT 0.998000 0.574000 1.059000 0.729000 ;
        RECT 0.544000 0.574000 1.059000 0.629000 ;
        END
    END SE
    PIN SI
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.655000 0.412000 0.790000 0.500000 ;
        RECT 0.655000 0.433000 0.838000 0.500000 ;
        END
    END SI
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 2.983000 1.078000 3.447000 1.280000 ;
        RECT 0.000000 1.120000 4.200000 1.280000 ;
        RECT 3.882000 1.078000 3.972000 1.280000 ;
        RECT 2.182000 1.078000 2.272000 1.280000 ;
        RECT 0.997000 1.065000 1.087000 1.280000 ;
        RECT 0.313000 1.078000 0.403000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 4.200000 0.080000 ;
        RECT 0.742000 -0.080000 0.833000 0.122000 ;
        RECT 4.057000 -0.080000 4.147000 0.211000 ;
        RECT 3.643000 -0.080000 3.733000 0.122000 ;
        RECT 2.286000 -0.080000 2.376000 0.308000 ;
        RECT 1.676000 -0.080000 1.766000 0.287000 ;
        RECT 0.231000 -0.080000 0.321000 0.409000 ;
        RECT 3.138000 -0.080000 3.199000 0.241000 ;
        RECT 0.231000 0.358000 0.329000 0.409000 ;
        END
    END VSS
    OBS
        LAYER Metal1 ;
        RECT 0.103000 0.719000 0.209000 0.913000 ;
        RECT 3.679000 0.931000 3.770000 1.040000 ;
        RECT 3.336000 0.277000 3.426000 0.412000 ;
        RECT 2.591000 0.576000 2.681000 0.752000 ;
        RECT 1.588000 0.926000 1.677000 1.019000 ;
        RECT 2.039000 0.150000 2.125000 0.344000 ;
        RECT 1.588000 0.933000 1.678000 1.019000 ;
        RECT 3.855000 0.348000 3.945000 0.429000 ;
        RECT 3.367000 0.917000 3.458000 0.998000 ;
        RECT 3.116000 0.800000 3.206000 0.881000 ;
        RECT 2.781000 0.807000 2.872000 0.888000 ;
        RECT 2.591000 0.917000 2.681000 0.998000 ;
        RECT 2.487000 0.262000 2.577000 0.343000 ;
        RECT 2.039000 0.263000 2.164000 0.344000 ;
        RECT 1.661000 0.514000 1.963000 0.595000 ;
        RECT 1.315000 0.193000 1.405000 0.274000 ;
        RECT 1.266000 0.769000 1.356000 0.850000 ;
        RECT 1.254000 0.329000 1.344000 0.410000 ;
        RECT 1.103000 0.179000 1.193000 0.260000 ;
        RECT 0.602000 0.724000 0.692000 0.805000 ;
        RECT 0.472000 0.343000 0.562000 0.424000 ;
        RECT 0.048000 0.319000 0.151000 0.400000 ;
        RECT 0.419000 0.700000 0.552000 0.779000 ;
        RECT 0.487000 0.302000 0.562000 0.424000 ;
        RECT 0.851000 0.302000 0.941000 0.373000 ;
        RECT 0.090000 0.719000 0.209000 0.788000 ;
        RECT 1.417000 0.926000 1.677000 0.988000 ;
        RECT 3.997000 0.374000 4.058000 0.986000 ;
        RECT 3.874000 0.544000 3.935000 0.876000 ;
        RECT 3.573000 0.357000 3.634000 0.876000 ;
        RECT 3.451000 0.467000 3.512000 0.745000 ;
        RECT 3.116000 0.800000 3.177000 0.998000 ;
        RECT 3.005000 0.152000 3.066000 0.412000 ;
        RECT 2.884000 0.262000 2.945000 0.521000 ;
        RECT 2.811000 0.690000 2.872000 0.888000 ;
        RECT 2.709000 0.152000 2.770000 0.289000 ;
        RECT 2.591000 0.454000 2.652000 0.752000 ;
        RECT 2.516000 0.262000 2.577000 0.399000 ;
        RECT 2.414000 0.807000 2.475000 0.888000 ;
        RECT 2.292000 0.698000 2.353000 1.008000 ;
        RECT 2.170000 0.563000 2.231000 0.899000 ;
        RECT 2.048000 0.563000 2.109000 0.706000 ;
        RECT 2.039000 0.150000 2.100000 0.618000 ;
        RECT 1.902000 0.226000 1.963000 0.899000 ;
        RECT 1.539000 0.368000 1.600000 0.857000 ;
        RECT 1.427000 0.219000 1.488000 0.423000 ;
        RECT 1.417000 0.619000 1.478000 0.988000 ;
        RECT 1.282000 0.329000 1.343000 0.674000 ;
        RECT 0.875000 0.933000 0.936000 1.050000 ;
        RECT 0.753000 0.795000 0.814000 0.936000 ;
        RECT 0.616000 0.154000 0.677000 0.248000 ;
        RECT 0.464000 0.858000 0.525000 1.050000 ;
        RECT 0.390000 0.369000 0.451000 0.755000 ;
        RECT 0.090000 0.319000 0.151000 0.788000 ;
        RECT 3.855000 0.374000 4.058000 0.429000 ;
        RECT 3.573000 0.821000 3.935000 0.876000 ;
        RECT 3.367000 0.931000 4.058000 0.986000 ;
        RECT 3.116000 0.800000 3.634000 0.855000 ;
        RECT 3.005000 0.357000 3.634000 0.412000 ;
        RECT 2.811000 0.690000 3.512000 0.745000 ;
        RECT 2.709000 0.152000 3.066000 0.207000 ;
        RECT 2.591000 0.943000 3.177000 0.998000 ;
        RECT 2.591000 0.576000 3.370000 0.631000 ;
        RECT 2.516000 0.344000 2.945000 0.399000 ;
        RECT 2.414000 0.807000 2.872000 0.862000 ;
        RECT 2.170000 0.563000 2.453000 0.618000 ;
        RECT 2.039000 0.563000 2.109000 0.618000 ;
        RECT 2.030000 0.150000 2.125000 0.205000 ;
        RECT 1.902000 0.844000 2.231000 0.899000 ;
        RECT 1.427000 0.368000 1.808000 0.423000 ;
        RECT 1.315000 0.219000 1.488000 0.274000 ;
        RECT 1.282000 0.619000 1.478000 0.674000 ;
        RECT 0.875000 0.933000 1.678000 0.988000 ;
        RECT 0.753000 0.795000 1.356000 0.850000 ;
        RECT 0.616000 0.193000 1.193000 0.248000 ;
        RECT 0.609000 0.881000 0.814000 0.936000 ;
        RECT 0.487000 0.302000 0.941000 0.357000 ;
        RECT 0.464000 0.995000 0.936000 1.050000 ;
        RECT 0.419000 0.724000 0.692000 0.779000 ;
        RECT 0.390000 0.700000 0.552000 0.755000 ;
        RECT 0.390000 0.369000 0.562000 0.424000 ;
        RECT 0.103000 0.858000 0.525000 0.913000 ;
        RECT 2.884000 0.467000 3.512000 0.521000 ;
        RECT 2.678000 0.235000 2.770000 0.289000 ;
        RECT 2.292000 0.698000 2.681000 0.752000 ;
        RECT 2.161000 0.454000 2.652000 0.508000 ;
        RECT 1.588000 0.954000 2.353000 1.008000 ;
        RECT 0.382000 0.154000 0.677000 0.208000 ;
        RECT 2.048000 0.150000 2.100000 0.706000 ;
        RECT 0.103000 0.319000 0.151000 0.913000 ;
        RECT 0.419000 0.369000 0.451000 0.779000 ;
    END
END SDFFHQX2

MACRO SDFFX2
    CLASS CORE ;
    FOREIGN SDFFX2 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 4.400000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER Metal1 ;
        RECT 0.213000 0.512000 0.329000 0.633000 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.057000 0.335000 1.191000 0.494000 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 3.696000 0.167000 3.787000 0.257000 ;
        RECT 3.589000 0.683000 3.680000 0.764000 ;
        RECT 3.589000 0.567000 3.659000 0.764000 ;
        RECT 3.557000 0.567000 3.659000 0.633000 ;
        RECT 3.540000 0.202000 3.601000 0.621000 ;
        RECT 3.540000 0.202000 3.787000 0.257000 ;
        RECT 3.540000 0.567000 3.659000 0.621000 ;
        RECT 3.557000 0.202000 3.589000 0.633000 ;
        RECT 3.589000 0.202000 3.601000 0.764000 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 4.085000 0.323000 4.167000 0.439000 ;
        RECT 4.059000 0.323000 4.167000 0.404000 ;
        RECT 4.000000 0.738000 4.091000 0.819000 ;
        RECT 4.105000 0.323000 4.167000 0.793000 ;
        RECT 4.000000 0.738000 4.167000 0.793000 ;
        END
    END QN
    PIN SE
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.020000 0.648000 1.111000 0.729000 ;
        RECT 0.547000 0.567000 0.667000 0.633000 ;
        RECT 1.020000 0.573000 1.081000 0.729000 ;
        RECT 1.019000 0.573000 1.081000 0.633000 ;
        RECT 0.547000 0.573000 1.081000 0.627000 ;
        END
    END SE
    PIN SI
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.672000 0.412000 0.765000 0.500000 ;
        RECT 0.672000 0.433000 0.843000 0.500000 ;
        END
    END SI
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 2.888000 1.078000 3.355000 1.280000 ;
        RECT 1.933000 1.078000 2.275000 1.280000 ;
        RECT 0.000000 1.120000 4.400000 1.280000 ;
        RECT 3.792000 1.078000 3.883000 1.280000 ;
        RECT 0.260000 1.078000 0.351000 1.280000 ;
        RECT 4.203000 1.078000 4.293000 1.280000 ;
        RECT 1.003000 1.065000 1.093000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 4.400000 0.080000 ;
        RECT 4.261000 -0.080000 4.352000 0.122000 ;
        RECT 3.909000 -0.080000 4.000000 0.122000 ;
        RECT 2.960000 -0.080000 3.051000 0.287000 ;
        RECT 1.685000 -0.080000 1.776000 0.287000 ;
        RECT 0.232000 -0.080000 0.323000 0.409000 ;
        RECT 3.483000 -0.080000 3.573000 0.122000 ;
        RECT 2.263000 -0.080000 2.353000 0.329000 ;
        RECT 0.747000 -0.080000 0.837000 0.122000 ;
        RECT 0.232000 0.358000 0.331000 0.409000 ;
        END
    END VSS
    OBS
        LAYER Metal1 ;
        RECT 3.944000 0.933000 4.035000 1.038000 ;
        RECT 3.589000 0.933000 3.680000 1.040000 ;
        RECT 3.173000 0.275000 3.264000 0.427000 ;
        RECT 2.560000 0.573000 2.651000 0.752000 ;
        RECT 2.536000 0.819000 2.627000 1.012000 ;
        RECT 1.587000 0.926000 1.677000 1.019000 ;
        RECT 1.587000 0.926000 1.679000 1.008000 ;
        RECT 3.696000 0.352000 3.787000 0.433000 ;
        RECT 3.275000 0.907000 3.365000 0.988000 ;
        RECT 3.021000 0.800000 3.112000 0.881000 ;
        RECT 2.619000 0.250000 2.709000 0.331000 ;
        RECT 2.179000 0.412000 2.269000 0.493000 ;
        RECT 2.055000 0.263000 2.156000 0.344000 ;
        RECT 2.035000 0.625000 2.125000 0.706000 ;
        RECT 1.660000 0.517000 1.953000 0.598000 ;
        RECT 1.323000 0.193000 1.413000 0.274000 ;
        RECT 1.263000 0.776000 1.353000 0.857000 ;
        RECT 1.261000 0.329000 1.352000 0.410000 ;
        RECT 1.109000 0.179000 1.200000 0.260000 ;
        RECT 0.605000 0.724000 0.696000 0.805000 ;
        RECT 0.475000 0.343000 0.565000 0.424000 ;
        RECT 0.048000 0.720000 0.152000 0.801000 ;
        RECT 0.048000 0.319000 0.152000 0.400000 ;
        RECT 3.133000 0.560000 3.224000 0.640000 ;
        RECT 2.376000 0.535000 2.467000 0.615000 ;
        RECT 0.424000 0.700000 0.555000 0.779000 ;
        RECT 3.036000 0.730000 3.112000 0.881000 ;
        RECT 0.489000 0.302000 0.565000 0.424000 ;
        RECT 0.856000 0.302000 0.947000 0.375000 ;
        RECT 3.753000 0.544000 3.815000 0.874000 ;
        RECT 3.021000 0.800000 3.083000 0.943000 ;
        RECT 2.205000 0.561000 2.267000 0.899000 ;
        RECT 1.537000 0.368000 1.599000 0.857000 ;
        RECT 1.415000 0.926000 1.679000 0.988000 ;
        RECT 0.757000 0.802000 0.819000 0.936000 ;
        RECT 3.876000 0.379000 3.937000 0.988000 ;
        RECT 3.464000 0.730000 3.525000 0.874000 ;
        RECT 3.303000 0.423000 3.364000 0.785000 ;
        RECT 3.203000 0.275000 3.264000 0.477000 ;
        RECT 2.811000 0.276000 2.872000 0.427000 ;
        RECT 2.560000 0.412000 2.621000 0.752000 ;
        RECT 2.331000 0.698000 2.392000 1.008000 ;
        RECT 2.055000 0.150000 2.116000 0.706000 ;
        RECT 1.895000 0.540000 1.956000 0.899000 ;
        RECT 1.892000 0.226000 1.953000 0.598000 ;
        RECT 1.435000 0.219000 1.496000 0.425000 ;
        RECT 1.415000 0.658000 1.476000 0.988000 ;
        RECT 1.291000 0.329000 1.352000 0.713000 ;
        RECT 0.880000 0.933000 0.941000 1.050000 ;
        RECT 0.620000 0.154000 0.681000 0.248000 ;
        RECT 0.467000 0.858000 0.528000 1.050000 ;
        RECT 0.424000 0.369000 0.485000 0.779000 ;
        RECT 0.091000 0.319000 0.152000 0.913000 ;
        RECT 1.895000 0.226000 1.953000 0.899000 ;
        RECT 1.660000 0.540000 1.956000 0.598000 ;
        RECT 1.435000 0.368000 1.599000 0.425000 ;
        RECT 3.464000 0.819000 3.815000 0.874000 ;
        RECT 3.275000 0.933000 4.035000 0.988000 ;
        RECT 3.036000 0.730000 3.525000 0.785000 ;
        RECT 2.619000 0.276000 2.872000 0.331000 ;
        RECT 2.536000 0.888000 3.083000 0.943000 ;
        RECT 2.179000 0.412000 2.621000 0.467000 ;
        RECT 2.020000 0.150000 2.116000 0.205000 ;
        RECT 1.895000 0.844000 2.267000 0.899000 ;
        RECT 1.435000 0.370000 1.819000 0.425000 ;
        RECT 1.323000 0.219000 1.496000 0.274000 ;
        RECT 1.291000 0.658000 1.476000 0.713000 ;
        RECT 0.880000 0.933000 1.679000 0.988000 ;
        RECT 0.757000 0.802000 1.353000 0.857000 ;
        RECT 0.620000 0.193000 1.200000 0.248000 ;
        RECT 0.612000 0.881000 0.819000 0.936000 ;
        RECT 0.489000 0.302000 0.947000 0.357000 ;
        RECT 0.467000 0.995000 0.941000 1.050000 ;
        RECT 0.424000 0.724000 0.696000 0.779000 ;
        RECT 0.424000 0.369000 0.565000 0.424000 ;
        RECT 0.091000 0.858000 0.528000 0.913000 ;
        RECT 3.696000 0.379000 3.937000 0.433000 ;
        RECT 3.203000 0.423000 3.364000 0.477000 ;
        RECT 2.811000 0.373000 3.264000 0.427000 ;
        RECT 2.627000 0.573000 3.224000 0.627000 ;
        RECT 2.560000 0.573000 3.112000 0.627000 ;
        RECT 2.331000 0.698000 2.651000 0.752000 ;
        RECT 2.205000 0.561000 2.467000 0.615000 ;
        RECT 1.587000 0.954000 2.392000 1.008000 ;
        RECT 0.384000 0.154000 0.681000 0.208000 ;
        RECT 3.036000 0.730000 3.083000 0.943000 ;
        RECT 0.475000 0.343000 0.485000 0.779000 ;
    END
END SDFFX2

MACRO OR4X4
    CLASS CORE ;
    FOREIGN OR4X4 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 2.000000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.683000 0.549000 0.882000 0.639000 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.405000 0.415000 0.592000 0.523000 ;
        RECT 0.937000 0.400000 1.030000 0.494000 ;
        RECT 0.499000 0.415000 0.592000 0.602000 ;
        RECT 0.405000 0.415000 1.030000 0.494000 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.299000 0.633000 0.401000 0.776000 ;
        RECT 0.303000 0.620000 0.397000 0.776000 ;
        RECT 1.128000 0.548000 1.222000 0.629000 ;
        RECT 0.934000 0.700000 1.207000 0.776000 ;
        RECT 0.299000 0.700000 0.423000 0.776000 ;
        RECT 1.143000 0.548000 1.207000 0.776000 ;
        RECT 0.299000 0.721000 1.207000 0.776000 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.220000 0.833000 0.424000 0.926000 ;
        RECT 1.178000 0.388000 1.271000 0.469000 ;
        RECT 0.129000 0.620000 0.193000 0.894000 ;
        RECT 1.302000 0.414000 1.365000 0.888000 ;
        RECT 0.129000 0.833000 0.424000 0.894000 ;
        RECT 1.178000 0.414000 1.365000 0.469000 ;
        RECT 0.129000 0.833000 1.365000 0.888000 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 2.000000 1.280000 ;
        RECT 1.394000 1.078000 1.488000 1.280000 ;
        RECT 1.791000 1.078000 1.884000 1.280000 ;
        RECT 0.050000 0.977000 0.143000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 2.000000 0.080000 ;
        RECT 1.292000 -0.080000 1.386000 0.122000 ;
        RECT 0.457000 -0.080000 0.551000 0.122000 ;
        RECT 1.769000 -0.080000 1.862000 0.122000 ;
        RECT 0.050000 -0.080000 0.143000 0.399000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.493000 0.344000 1.675000 0.793000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 0.713000 0.154000 0.807000 0.346000 ;
        RECT 0.248000 0.221000 0.342000 0.414000 ;
        RECT 1.758000 0.500000 1.851000 0.581000 ;
        RECT 0.711000 0.944000 0.804000 1.025000 ;
        RECT 1.773000 0.223000 1.836000 0.999000 ;
        RECT 0.566000 0.223000 0.629000 0.345000 ;
        RECT 0.711000 0.944000 1.836000 0.999000 ;
        RECT 0.248000 0.290000 0.629000 0.345000 ;
        RECT 0.566000 0.223000 1.836000 0.277000 ;
    END
END OR4X4

MACRO OR4X2
    CLASS CORE ;
    FOREIGN OR4X2 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 1.100000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.039000 0.433000 0.151000 0.567000 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.222000 0.167000 0.364000 0.264000 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.406000 0.527000 0.556000 0.633000 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.664000 0.700000 0.878000 0.767000 ;
        RECT 0.664000 0.552000 0.728000 0.767000 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 1.100000 1.280000 ;
        RECT 0.742000 1.078000 0.836000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 1.100000 0.080000 ;
        RECT 0.551000 -0.080000 0.646000 0.122000 ;
        RECT 0.050000 -0.080000 0.144000 0.122000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.942000 0.182000 1.061000 0.375000 ;
        RECT 0.953000 0.700000 1.061000 1.010000 ;
        RECT 0.997000 0.182000 1.061000 1.010000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 0.812000 0.462000 0.918000 0.576000 ;
        RECT 0.050000 0.731000 0.144000 0.924000 ;
        RECT 0.575000 0.320000 0.669000 0.401000 ;
        RECT 0.215000 0.320000 0.285000 0.388000 ;
        RECT 0.812000 0.333000 0.876000 0.576000 ;
        RECT 0.215000 0.320000 0.279000 0.717000 ;
        RECT 0.081000 0.662000 0.144000 0.924000 ;
        RECT 0.285000 0.333000 0.876000 0.388000 ;
        RECT 0.081000 0.662000 0.279000 0.717000 ;
    END
END OR4X2

MACRO OR3X4
    CLASS CORE ;
    FOREIGN OR3X4 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 1.600000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.392000 0.567000 0.548000 0.694000 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.667000 0.457000 0.758000 0.583000 ;
        RECT 0.172000 0.431000 0.264000 0.512000 ;
        RECT 0.172000 0.439000 0.298000 0.512000 ;
        RECT 0.172000 0.457000 0.758000 0.512000 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.038000 0.681000 0.215000 0.775000 ;
        RECT 0.124000 0.604000 0.215000 0.775000 ;
        RECT 0.154000 0.700000 0.236000 0.804000 ;
        RECT 0.038000 0.700000 0.236000 0.775000 ;
        RECT 0.634000 0.704000 0.769000 0.767000 ;
        RECT 0.855000 0.413000 0.917000 0.758000 ;
        RECT 0.634000 0.704000 0.696000 0.804000 ;
        RECT 0.154000 0.604000 0.215000 0.804000 ;
        RECT 0.831000 0.700000 0.917000 0.758000 ;
        RECT 0.855000 0.413000 0.966000 0.468000 ;
        RECT 0.154000 0.749000 0.696000 0.804000 ;
        RECT 0.634000 0.704000 0.917000 0.758000 ;
        END
    END C
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 1.600000 1.280000 ;
        RECT 1.418000 0.983000 1.510000 1.280000 ;
        RECT 1.061000 0.983000 1.153000 1.280000 ;
        RECT 0.048000 1.078000 0.140000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 1.600000 0.080000 ;
        RECT 1.403000 -0.080000 1.495000 0.122000 ;
        RECT 0.529000 -0.080000 0.621000 0.222000 ;
        RECT 0.958000 -0.080000 1.049000 0.122000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.104000 0.331000 1.207000 0.767000 ;
        RECT 1.104000 0.679000 1.339000 0.767000 ;
        RECT 1.104000 0.331000 1.274000 0.412000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 0.739000 0.213000 0.835000 0.358000 ;
        RECT 0.739000 0.162000 0.831000 0.358000 ;
        RECT 0.322000 0.162000 0.413000 0.358000 ;
        RECT 1.332000 0.532000 1.463000 0.613000 ;
        RECT 0.555000 0.896000 0.646000 0.977000 ;
        RECT 1.401000 0.213000 1.463000 0.898000 ;
        RECT 0.791000 0.843000 0.853000 0.951000 ;
        RECT 0.835000 0.213000 1.463000 0.268000 ;
        RECT 0.791000 0.843000 1.463000 0.898000 ;
        RECT 0.739000 0.213000 1.332000 0.268000 ;
        RECT 0.555000 0.896000 0.853000 0.951000 ;
        RECT 0.322000 0.304000 0.835000 0.358000 ;
    END
END OR3X4

MACRO OR3X2
    CLASS CORE ;
    FOREIGN OR3X2 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 1.100000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.186000 0.567000 0.322000 0.668000 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.411000 0.423000 0.506000 0.518000 ;
        RECT 0.383000 0.423000 0.539000 0.507000 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.586000 0.601000 0.700000 0.775000 ;
        END
    END C
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 1.100000 1.280000 ;
        RECT 0.722000 1.078000 0.817000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 1.100000 0.080000 ;
        RECT 0.744000 -0.080000 0.839000 0.211000 ;
        RECT 0.281000 -0.080000 0.375000 0.122000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.944000 0.182000 1.061000 0.375000 ;
        RECT 0.956000 0.182000 1.061000 0.500000 ;
        RECT 0.944000 0.705000 1.039000 1.010000 ;
        RECT 0.975000 0.182000 1.039000 1.010000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 0.161000 0.756000 0.256000 0.949000 ;
        RECT 0.046000 0.300000 0.147000 0.381000 ;
        RECT 0.787000 0.481000 0.862000 0.568000 ;
        RECT 0.787000 0.313000 0.851000 0.568000 ;
        RECT 0.046000 0.300000 0.110000 0.811000 ;
        RECT 0.161000 0.313000 0.851000 0.368000 ;
        RECT 0.147000 0.313000 0.787000 0.368000 ;
        RECT 0.046000 0.756000 0.256000 0.811000 ;
        RECT 0.046000 0.313000 0.256000 0.368000 ;
    END
END OR3X2

MACRO OR2X4
    CLASS CORE ;
    FOREIGN OR2X4 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 1.100000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.039000 0.392000 0.144000 0.556000 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.343000 0.479000 0.511000 0.663000 ;
        END
    END B
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 1.100000 1.280000 ;
        RECT 0.794000 1.078000 0.889000 1.280000 ;
        RECT 0.417000 1.078000 0.511000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 1.100000 0.080000 ;
        RECT 0.461000 -0.080000 0.556000 0.214000 ;
        RECT 0.828000 -0.080000 0.922000 0.122000 ;
        RECT 0.050000 -0.080000 0.144000 0.290000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.589000 0.300000 0.694000 0.633000 ;
        RECT 0.606000 0.624000 0.696000 0.733000 ;
        RECT 0.606000 0.300000 0.694000 0.733000 ;
        RECT 0.606000 0.652000 0.700000 0.733000 ;
        RECT 0.589000 0.324000 0.733000 0.405000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 0.772000 0.500000 0.867000 0.581000 ;
        RECT 0.214000 0.276000 0.344000 0.357000 ;
        RECT 0.050000 0.669000 0.278000 0.750000 ;
        RECT 0.772000 0.500000 0.836000 0.843000 ;
        RECT 0.214000 0.276000 0.278000 0.843000 ;
        RECT 0.214000 0.788000 0.836000 0.843000 ;
    END
END OR2X4

MACRO OR2X2
    CLASS CORE ;
    FOREIGN OR2X2 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 0.700000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.037000 0.393000 0.138000 0.544000 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.212000 0.414000 0.337000 0.558000 ;
        END
    END B
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 0.700000 1.280000 ;
        RECT 0.345000 1.078000 0.435000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 0.700000 0.080000 ;
        RECT 0.345000 -0.080000 0.435000 0.122000 ;
        RECT 0.048000 -0.080000 0.138000 0.122000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.546000 0.721000 0.650000 0.914000 ;
        RECT 0.548000 0.196000 0.650000 0.389000 ;
        RECT 0.589000 0.196000 0.650000 0.914000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 0.399000 0.502000 0.528000 0.583000 ;
        RECT 0.196000 0.252000 0.286000 0.333000 ;
        RECT 0.048000 0.721000 0.138000 0.802000 ;
        RECT 0.399000 0.279000 0.460000 0.776000 ;
        RECT 0.048000 0.721000 0.460000 0.776000 ;
        RECT 0.196000 0.279000 0.460000 0.333000 ;
    END
END OR2X2

MACRO OAI33X2
    CLASS CORE ;
    FOREIGN OAI33X2 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 2.300000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.473000 0.567000 1.659000 0.651000 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.285000 0.439000 1.358000 0.512000 ;
        RECT 1.285000 0.439000 1.347000 0.555000 ;
        RECT 1.779000 0.457000 1.840000 0.555000 ;
        RECT 1.285000 0.457000 1.840000 0.512000 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.091000 0.300000 1.182000 0.455000 ;
        RECT 1.993000 0.567000 2.055000 0.761000 ;
        RECT 1.119000 0.300000 1.181000 0.761000 ;
        RECT 1.119000 0.706000 2.055000 0.761000 ;
        END
    END A2
    PIN B0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.477000 0.549000 0.670000 0.633000 ;
        END
    END B0
    PIN B1
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.765000 0.433000 0.877000 0.556000 ;
        RECT 0.765000 0.433000 0.862000 0.627000 ;
        RECT 0.294000 0.433000 0.383000 0.556000 ;
        RECT 0.292000 0.475000 0.383000 0.556000 ;
        RECT 0.294000 0.433000 0.877000 0.488000 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.058000 0.536000 0.139000 0.627000 ;
        RECT 0.051000 0.536000 0.142000 0.617000 ;
        RECT 0.965000 0.535000 1.056000 0.615000 ;
        RECT 0.965000 0.535000 1.027000 0.748000 ;
        RECT 0.078000 0.536000 0.139000 0.748000 ;
        RECT 0.078000 0.693000 1.027000 0.748000 ;
        END
    END B2
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 2.300000 1.280000 ;
        RECT 2.053000 1.078000 2.145000 1.280000 ;
        RECT 1.045000 1.078000 1.137000 1.280000 ;
        RECT 0.048000 0.817000 0.139000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 2.300000 0.080000 ;
        RECT 0.544000 -0.080000 0.635000 0.211000 ;
        RECT 0.048000 -0.080000 0.139000 0.211000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.549000 0.839000 1.641000 1.050000 ;
        RECT 0.541000 0.826000 0.633000 0.907000 ;
        RECT 2.116000 0.324000 2.178000 0.894000 ;
        RECT 2.065000 0.833000 2.178000 0.894000 ;
        RECT 1.264000 0.324000 2.178000 0.379000 ;
        RECT 0.541000 0.839000 2.178000 0.894000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 0.842000 0.158000 0.903000 0.379000 ;
        RECT 0.842000 0.158000 2.090000 0.213000 ;
        RECT 0.260000 0.324000 0.903000 0.379000 ;
    END
END OAI33X2

MACRO OAI32X2
    CLASS CORE ;
    FOREIGN OAI32X2 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 2.000000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.463000 0.614000 0.584000 0.761000 ;
        RECT 0.423000 0.706000 0.584000 0.761000 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.766000 0.492000 0.871000 0.631000 ;
        RECT 0.777000 0.479000 0.871000 0.631000 ;
        RECT 0.302000 0.479000 0.395000 0.560000 ;
        RECT 0.302000 0.492000 0.871000 0.546000 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.116000 0.613000 0.209000 0.706000 ;
        RECT 0.961000 0.614000 1.055000 0.706000 ;
        RECT 0.116000 0.573000 0.194000 0.706000 ;
        RECT 0.116000 0.639000 0.337000 0.706000 ;
        RECT 0.961000 0.614000 1.025000 0.771000 ;
        RECT 0.712000 0.717000 0.775000 0.887000 ;
        RECT 0.274000 0.639000 0.337000 0.887000 ;
        RECT 0.274000 0.832000 0.775000 0.887000 ;
        RECT 0.712000 0.717000 1.025000 0.771000 ;
        RECT 0.059000 0.573000 0.194000 0.627000 ;
        END
    END A2
    PIN B0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.322000 0.598000 1.467000 0.761000 ;
        END
    END B0
    PIN B1
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.150000 0.479000 1.245000 0.623000 ;
        RECT 1.558000 0.479000 1.652000 0.560000 ;
        RECT 1.150000 0.479000 1.213000 0.627000 ;
        RECT 1.150000 0.479000 1.652000 0.533000 ;
        END
    END B1
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 2.000000 1.280000 ;
        RECT 1.803000 1.078000 1.897000 1.280000 ;
        RECT 1.076000 1.078000 1.169000 1.280000 ;
        RECT 0.050000 0.877000 0.143000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 2.000000 0.080000 ;
        RECT 0.603000 -0.080000 0.697000 0.211000 ;
        RECT 0.094000 -0.080000 0.187000 0.211000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.675000 0.839000 1.822000 0.964000 ;
        RECT 1.532000 0.343000 1.625000 0.424000 ;
        RECT 1.439000 0.896000 1.533000 0.977000 ;
        RECT 1.077000 0.343000 1.171000 0.424000 ;
        RECT 0.556000 0.969000 0.650000 1.050000 ;
        RECT 0.850000 0.967000 0.983000 1.037000 ;
        RECT 1.532000 0.343000 1.696000 0.411000 ;
        RECT 1.759000 0.356000 1.822000 0.964000 ;
        RECT 0.920000 0.910000 0.983000 1.037000 ;
        RECT 1.077000 0.356000 1.822000 0.411000 ;
        RECT 0.556000 0.982000 0.983000 1.037000 ;
        RECT 0.920000 0.910000 1.822000 0.964000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 1.227000 0.150000 1.450000 0.231000 ;
        RECT 0.837000 0.343000 0.931000 0.424000 ;
        RECT 0.270000 0.343000 0.493000 0.424000 ;
        RECT 0.868000 0.163000 0.931000 0.424000 ;
        RECT 0.868000 0.163000 1.450000 0.218000 ;
        RECT 0.493000 0.356000 0.837000 0.411000 ;
    END
END OAI32X2

MACRO OAI31X2
    CLASS CORE ;
    FOREIGN OAI31X2 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 1.600000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.479000 0.567000 0.673000 0.668000 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.811000 0.539000 0.902000 0.620000 ;
        RECT 0.294000 0.539000 0.393000 0.620000 ;
        RECT 0.811000 0.445000 0.873000 0.620000 ;
        RECT 0.331000 0.445000 0.393000 0.620000 ;
        RECT 0.413000 0.439000 0.475000 0.500000 ;
        RECT 0.331000 0.445000 0.873000 0.500000 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.143000 0.700000 0.236000 0.792000 ;
        RECT 0.947000 0.706000 1.037000 0.792000 ;
        RECT 0.991000 0.614000 1.083000 0.695000 ;
        RECT 0.113000 0.614000 0.205000 0.695000 ;
        RECT 0.975000 0.627000 1.083000 0.695000 ;
        RECT 0.975000 0.627000 1.037000 0.792000 ;
        RECT 0.143000 0.614000 0.205000 0.792000 ;
        RECT 0.143000 0.737000 1.037000 0.792000 ;
        RECT 0.991000 0.614000 1.037000 0.792000 ;
        END
    END A2
    PIN B0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.282000 0.567000 1.399000 0.719000 ;
        END
    END B0
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 1.600000 1.280000 ;
        RECT 1.445000 0.821000 1.537000 1.280000 ;
        RECT 0.048000 0.877000 0.140000 1.280000 ;
        RECT 1.067000 1.078000 1.158000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 1.600000 0.080000 ;
        RECT 0.932000 -0.080000 1.024000 0.122000 ;
        RECT 0.199000 -0.080000 0.291000 0.122000 ;
        RECT 0.555000 -0.080000 0.646000 0.122000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.154000 0.804000 1.343000 0.911000 ;
        RECT 0.544000 0.856000 0.636000 1.049000 ;
        RECT 1.277000 0.343000 1.368000 0.439000 ;
        RECT 1.125000 0.839000 1.343000 0.911000 ;
        RECT 1.277000 0.343000 1.339000 0.512000 ;
        RECT 1.154000 0.457000 1.216000 0.911000 ;
        RECT 1.154000 0.457000 1.339000 0.512000 ;
        RECT 0.544000 0.856000 1.343000 0.911000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 0.711000 0.151000 0.859000 0.365000 ;
        RECT 0.404000 0.298000 0.496000 0.379000 ;
        RECT 0.048000 0.298000 0.140000 0.379000 ;
        RECT 0.797000 0.151000 0.859000 0.390000 ;
        RECT 0.048000 0.324000 0.496000 0.379000 ;
        RECT 0.797000 0.336000 1.174000 0.390000 ;
        RECT 0.404000 0.311000 0.711000 0.365000 ;
    END
END OAI31X2

MACRO OAI2BB1X4
    CLASS CORE ;
    FOREIGN OAI2BB1X4 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 1.800000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A0N
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.331000 0.539000 0.502000 0.633000 ;
        END
    END A0N
    PIN A1N
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.038000 0.481000 0.142000 0.633000 ;
        END
    END A1N
    PIN B0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.578000 0.539000 0.824000 0.633000 ;
        END
    END B0
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 1.800000 1.280000 ;
        RECT 1.190000 0.877000 1.283000 1.280000 ;
        RECT 0.841000 0.877000 0.934000 1.280000 ;
        RECT 0.049000 0.747000 0.142000 1.280000 ;
        RECT 0.475000 0.944000 0.567000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 1.800000 0.080000 ;
        RECT 0.747000 -0.080000 0.840000 0.212000 ;
        RECT 0.398000 -0.080000 0.491000 0.212000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.478000 0.567000 1.582000 0.900000 ;
        RECT 1.561000 0.170000 1.669000 0.251000 ;
        RECT 1.216000 0.170000 1.309000 0.251000 ;
        RECT 1.016000 0.688000 1.139000 0.769000 ;
        RECT 0.667000 0.688000 0.760000 0.769000 ;
        RECT 1.557000 0.183000 1.669000 0.251000 ;
        RECT 1.216000 0.170000 1.320000 0.238000 ;
        RECT 0.667000 0.701000 0.779000 0.769000 ;
        RECT 1.557000 0.183000 1.620000 0.621000 ;
        RECT 1.561000 0.170000 1.620000 0.621000 ;
        RECT 1.216000 0.183000 1.669000 0.238000 ;
        RECT 0.667000 0.701000 1.582000 0.756000 ;
        RECT 1.478000 0.567000 1.620000 0.621000 ;
        RECT 1.561000 0.170000 1.582000 0.900000 ;
        RECT 1.557000 0.183000 1.561000 0.900000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 1.402000 0.319000 1.495000 0.424000 ;
        RECT 0.256000 0.732000 0.349000 1.037000 ;
        RECT 0.049000 0.151000 0.142000 0.344000 ;
        RECT 0.955000 0.280000 1.047000 0.374000 ;
        RECT 1.065000 0.525000 1.414000 0.606000 ;
        RECT 0.910000 0.430000 0.972000 0.580000 ;
        RECT 0.205000 0.289000 0.267000 0.788000 ;
        RECT 0.588000 0.319000 0.650000 0.375000 ;
        RECT 0.205000 0.732000 0.349000 0.788000 ;
        RECT 0.910000 0.525000 1.414000 0.580000 ;
        RECT 0.588000 0.319000 1.495000 0.374000 ;
        RECT 0.573000 0.320000 0.650000 0.375000 ;
        RECT 0.349000 0.430000 0.972000 0.485000 ;
        RECT 0.267000 0.430000 0.910000 0.485000 ;
        RECT 0.205000 0.430000 0.650000 0.485000 ;
        RECT 0.049000 0.289000 0.267000 0.344000 ;
        RECT 0.573000 0.320000 1.495000 0.374000 ;
        RECT 0.256000 0.289000 0.267000 1.037000 ;
    END
END OAI2BB1X4

MACRO OAI2BB1X2
    CLASS CORE ;
    FOREIGN OAI2BB1X2 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 1.300000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A0N
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.359000 0.567000 0.568000 0.633000 ;
        RECT 0.359000 0.542000 0.423000 0.633000 ;
        END
    END A0N
    PIN A1N
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.060000 0.400000 0.165000 0.533000 ;
        END
    END A1N
    PIN B0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.535000 0.379000 0.703000 0.507000 ;
        END
    END B0
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 1.300000 1.280000 ;
        RECT 1.013000 1.078000 1.109000 1.280000 ;
        RECT 0.642000 0.972000 0.737000 1.280000 ;
        RECT 0.203000 1.078000 0.298000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 1.300000 0.080000 ;
        RECT 0.422000 -0.080000 0.518000 0.289000 ;
        RECT 1.154000 -0.080000 1.249000 0.289000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.822000 0.676000 0.917000 0.757000 ;
        RECT 0.794000 0.265000 0.889000 0.346000 ;
        RECT 0.989000 0.292000 1.054000 0.627000 ;
        RECT 0.968000 0.573000 1.033000 0.731000 ;
        RECT 0.822000 0.676000 1.033000 0.731000 ;
        RECT 0.968000 0.573000 1.054000 0.627000 ;
        RECT 0.794000 0.292000 1.054000 0.346000 ;
        RECT 0.989000 0.292000 1.033000 0.731000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 0.768000 0.468000 0.864000 0.549000 ;
        RECT 0.428000 0.768000 0.523000 0.849000 ;
        RECT 0.051000 0.254000 0.146000 0.335000 ;
        RECT 0.768000 0.468000 0.833000 0.621000 ;
        RECT 0.691000 0.567000 0.756000 0.823000 ;
        RECT 0.229000 0.280000 0.294000 0.823000 ;
        RECT 0.229000 0.768000 0.756000 0.823000 ;
        RECT 0.051000 0.280000 0.294000 0.335000 ;
        RECT 0.691000 0.567000 0.833000 0.621000 ;
    END
END OAI2BB1X2

MACRO OAI22X2
    CLASS CORE ;
    FOREIGN OAI22X2 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 1.600000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.843000 0.560000 0.948000 0.664000 ;
        RECT 0.843000 0.573000 1.009000 0.664000 ;
        RECT 1.343000 0.583000 1.434000 0.664000 ;
        RECT 0.843000 0.610000 1.434000 0.664000 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.104000 0.412000 1.239000 0.554000 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.048000 0.398000 0.140000 0.554000 ;
        RECT 0.663000 0.473000 0.754000 0.554000 ;
        RECT 0.661000 0.473000 0.754000 0.540000 ;
        RECT 0.661000 0.398000 0.723000 0.540000 ;
        RECT 0.663000 0.398000 0.723000 0.554000 ;
        RECT 0.048000 0.398000 0.723000 0.452000 ;
        END
    END B0
    PIN B1
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.339000 0.508000 0.558000 0.589000 ;
        RECT 0.236000 0.535000 0.298000 0.627000 ;
        RECT 0.236000 0.535000 0.558000 0.589000 ;
        END
    END B1
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 1.600000 1.280000 ;
        RECT 1.096000 0.911000 1.188000 1.280000 ;
        RECT 0.404000 0.911000 0.496000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 1.600000 0.080000 ;
        RECT 0.070000 -0.080000 0.162000 0.122000 ;
        RECT 0.555000 -0.080000 0.646000 0.122000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.441000 0.720000 1.558000 0.833000 ;
        RECT 1.282000 0.746000 1.558000 0.833000 ;
        RECT 1.282000 0.746000 1.364000 0.894000 ;
        RECT 1.309000 0.262000 1.401000 0.343000 ;
        RECT 0.954000 0.262000 1.045000 0.343000 ;
        RECT 0.752000 0.720000 0.843000 0.801000 ;
        RECT 0.048000 0.720000 0.140000 0.801000 ;
        RECT 1.496000 0.288000 1.558000 0.833000 ;
        RECT 0.954000 0.288000 1.558000 0.343000 ;
        RECT 0.048000 0.746000 1.558000 0.801000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 0.760000 0.261000 0.851000 0.342000 ;
        RECT 0.404000 0.261000 0.496000 0.342000 ;
        RECT 0.048000 0.261000 0.140000 0.342000 ;
        RECT 0.048000 0.287000 0.851000 0.342000 ;
    END
END OAI22X2

MACRO OAI222X2
    CLASS CORE ;
    FOREIGN OAI222X2 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 2.600000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.208000 0.662000 1.297000 0.767000 ;
        RECT 1.129000 0.700000 1.341000 0.767000 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.961000 0.560000 1.051000 0.640000 ;
        RECT 0.990000 0.552000 1.051000 0.640000 ;
        RECT 1.362000 0.552000 1.422000 0.617000 ;
        RECT 1.362000 0.562000 1.535000 0.617000 ;
        RECT 0.990000 0.552000 1.422000 0.607000 ;
        RECT 0.923000 0.573000 1.051000 0.627000 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.436000 0.662000 0.651000 0.743000 ;
        RECT 0.576000 0.662000 0.637000 0.761000 ;
        END
    END B0
    PIN B1
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.152000 0.546000 0.242000 0.627000 ;
        RECT 0.152000 0.552000 0.290000 0.627000 ;
        RECT 0.152000 0.552000 0.827000 0.607000 ;
        END
    END B1
    PIN C0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.943000 0.498000 2.043000 0.633000 ;
        END
    END C0
    PIN C1
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 2.125000 0.675000 2.185000 0.743000 ;
        RECT 1.673000 0.573000 1.733000 0.743000 ;
        RECT 2.125000 0.675000 2.214000 0.730000 ;
        RECT 1.673000 0.688000 2.185000 0.743000 ;
        RECT 1.616000 0.573000 1.733000 0.627000 ;
        END
    END C1
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 2.600000 1.280000 ;
        RECT 2.190000 0.984000 2.280000 1.280000 ;
        RECT 1.507000 0.984000 1.597000 1.280000 ;
        RECT 0.835000 0.984000 0.924000 1.280000 ;
        RECT 0.163000 0.984000 0.252000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 2.600000 0.080000 ;
        RECT 0.383000 -0.080000 0.473000 0.211000 ;
        RECT 0.047000 -0.080000 0.137000 0.211000 ;
        RECT 0.762000 -0.080000 0.851000 0.211000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.849000 0.839000 1.964000 0.920000 ;
        RECT 1.154000 0.839000 1.271000 0.920000 ;
        RECT 0.499000 0.839000 0.588000 0.920000 ;
        RECT 2.274000 0.331000 2.335000 0.888000 ;
        RECT 2.136000 0.833000 2.197000 0.894000 ;
        RECT 2.136000 0.833000 2.335000 0.888000 ;
        RECT 1.861000 0.331000 2.335000 0.386000 ;
        RECT 0.499000 0.839000 2.197000 0.894000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 1.114000 0.302000 1.203000 0.399000 ;
        RECT 0.573000 0.212000 0.662000 0.357000 ;
        RECT 0.215000 0.318000 0.305000 0.399000 ;
        RECT 1.686000 0.158000 1.746000 0.327000 ;
        RECT 0.573000 0.212000 0.633000 0.373000 ;
        RECT 1.686000 0.193000 2.487000 0.248000 ;
        RECT 0.945000 0.158000 1.746000 0.213000 ;
        RECT 0.573000 0.302000 1.572000 0.357000 ;
        RECT 0.215000 0.318000 0.633000 0.373000 ;
    END
END OAI222X2

MACRO OAI221X2
    CLASS CORE ;
    FOREIGN OAI221X2 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 2.300000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.104000 0.662000 1.196000 0.767000 ;
        RECT 1.024000 0.700000 1.240000 0.767000 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.863000 0.560000 0.954000 0.640000 ;
        RECT 0.863000 0.560000 1.004000 0.627000 ;
        RECT 1.257000 0.552000 1.319000 0.617000 ;
        RECT 0.942000 0.552000 1.004000 0.627000 ;
        RECT 1.257000 0.562000 1.512000 0.617000 ;
        RECT 0.942000 0.552000 1.319000 0.607000 ;
        RECT 0.942000 0.552000 0.954000 0.640000 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.327000 0.662000 0.547000 0.743000 ;
        RECT 0.411000 0.662000 0.473000 0.761000 ;
        END
    END B0
    PIN B1
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.113000 0.546000 0.204000 0.627000 ;
        RECT 0.113000 0.552000 0.740000 0.607000 ;
        RECT 0.058000 0.573000 0.204000 0.627000 ;
        END
    END B1
    PIN C0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.647000 0.567000 1.903000 0.633000 ;
        END
    END C0
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 2.300000 1.280000 ;
        RECT 1.817000 0.900000 1.909000 1.280000 ;
        RECT 0.734000 0.984000 0.826000 1.280000 ;
        RECT 1.421000 0.984000 1.512000 1.280000 ;
        RECT 0.048000 0.929000 0.139000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 2.300000 0.080000 ;
        RECT 0.777000 -0.080000 0.869000 0.211000 ;
        RECT 0.391000 -0.080000 0.483000 0.211000 ;
        RECT 0.048000 -0.080000 0.139000 0.211000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.914000 0.345000 2.032000 0.440000 ;
        RECT 1.624000 0.823000 1.716000 0.904000 ;
        RECT 1.078000 0.839000 1.169000 0.920000 ;
        RECT 0.391000 0.839000 0.483000 0.920000 ;
        RECT 1.654000 0.775000 1.732000 0.839000 ;
        RECT 1.970000 0.345000 2.032000 0.830000 ;
        RECT 1.914000 0.318000 1.976000 0.440000 ;
        RECT 1.654000 0.775000 1.716000 0.904000 ;
        RECT 1.003000 0.839000 1.169000 0.900000 ;
        RECT 1.654000 0.775000 2.032000 0.830000 ;
        RECT 0.391000 0.839000 1.716000 0.894000 ;
        RECT 1.970000 0.318000 1.976000 0.830000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 0.584000 0.217000 0.676000 0.357000 ;
        RECT 1.137000 0.302000 1.228000 0.399000 ;
        RECT 0.220000 0.318000 0.311000 0.399000 ;
        RECT 1.721000 0.158000 1.783000 0.327000 ;
        RECT 0.584000 0.217000 0.646000 0.373000 ;
        RECT 1.721000 0.193000 2.162000 0.248000 ;
        RECT 0.965000 0.158000 1.783000 0.213000 ;
        RECT 0.584000 0.302000 1.604000 0.357000 ;
        RECT 0.220000 0.318000 0.646000 0.373000 ;
    END
END OAI221X2

MACRO OAI21X4
    CLASS CORE ;
    FOREIGN OAI21X4 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 2.000000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.028000 0.505000 1.121000 0.586000 ;
        RECT 0.336000 0.533000 0.584000 0.614000 ;
        RECT 0.423000 0.533000 0.492000 0.627000 ;
        RECT 1.028000 0.440000 1.091000 0.586000 ;
        RECT 0.521000 0.440000 0.584000 0.614000 ;
        RECT 0.521000 0.440000 1.091000 0.495000 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.116000 0.533000 0.209000 0.627000 ;
        RECT 0.689000 0.550000 0.788000 0.633000 ;
        RECT 0.131000 0.533000 0.209000 0.633000 ;
        RECT 0.689000 0.550000 0.752000 0.743000 ;
        RECT 0.146000 0.533000 0.209000 0.743000 ;
        RECT 0.689000 0.550000 0.937000 0.605000 ;
        RECT 0.146000 0.688000 0.752000 0.743000 ;
        RECT 0.059000 0.573000 0.209000 0.627000 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.262000 0.560000 1.488000 0.640000 ;
        END
    END B0
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 2.000000 1.280000 ;
        RECT 0.766000 0.947000 0.860000 1.280000 ;
        RECT 1.660000 0.883000 1.753000 1.280000 ;
        RECT 1.306000 0.883000 1.399000 1.280000 ;
        RECT 0.050000 0.847000 0.143000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 2.000000 0.080000 ;
        RECT 0.953000 -0.080000 1.047000 0.211000 ;
        RECT 0.248000 -0.080000 0.342000 0.211000 ;
        RECT 0.601000 -0.080000 0.694000 0.211000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.675000 0.331000 1.809000 0.440000 ;
        RECT 1.675000 0.331000 1.780000 0.767000 ;
        RECT 1.715000 0.313000 1.809000 0.440000 ;
        RECT 1.482000 0.695000 1.576000 0.776000 ;
        RECT 1.129000 0.695000 1.223000 0.776000 ;
        RECT 0.402000 0.798000 0.496000 0.879000 ;
        RECT 1.715000 0.313000 1.780000 0.767000 ;
        RECT 1.129000 0.695000 1.193000 0.865000 ;
        RECT 1.329000 0.331000 1.809000 0.386000 ;
        RECT 1.129000 0.708000 1.780000 0.763000 ;
        RECT 0.402000 0.811000 1.193000 0.865000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 1.506000 0.150000 1.599000 0.231000 ;
        RECT 1.153000 0.150000 1.247000 0.231000 ;
        RECT 0.050000 0.226000 0.143000 0.307000 ;
        RECT 1.153000 0.150000 1.216000 0.386000 ;
        RECT 0.080000 0.226000 0.143000 0.386000 ;
        RECT 1.247000 0.163000 1.506000 0.218000 ;
        RECT 0.080000 0.331000 1.216000 0.386000 ;
    END
END OAI21X4

MACRO OAI21X2
    CLASS CORE ;
    FOREIGN OAI21X2 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 1.400000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.650000 0.605000 0.740000 0.686000 ;
        RECT 0.119000 0.433000 0.232000 0.514000 ;
        RECT 0.118000 0.439000 0.232000 0.514000 ;
        RECT 0.650000 0.460000 0.711000 0.686000 ;
        RECT 0.057000 0.439000 0.232000 0.494000 ;
        RECT 0.118000 0.460000 0.711000 0.514000 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.323000 0.614000 0.488000 0.707000 ;
        RECT 0.323000 0.614000 0.562000 0.695000 ;
        RECT 0.407000 0.614000 0.473000 0.761000 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.875000 0.551000 1.179000 0.632000 ;
        END
    END B0
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 1.400000 1.280000 ;
        RECT 0.949000 1.078000 1.039000 1.280000 ;
        RECT 0.398000 1.078000 0.488000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 1.400000 0.080000 ;
        RECT 0.642000 -0.080000 0.732000 0.280000 ;
        RECT 0.249000 -0.080000 0.339000 0.122000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.151000 0.865000 1.283000 0.946000 ;
        RECT 1.023000 0.263000 1.114000 0.344000 ;
        RECT 0.748000 0.865000 0.838000 0.946000 ;
        RECT 0.048000 0.865000 0.138000 0.946000 ;
        RECT 1.282000 0.311000 1.343000 0.920000 ;
        RECT 1.053000 0.263000 1.114000 0.365000 ;
        RECT 0.048000 0.865000 1.343000 0.920000 ;
        RECT 1.053000 0.311000 1.343000 0.365000 ;
        RECT 1.282000 0.311000 1.283000 0.946000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 1.214000 0.175000 1.305000 0.256000 ;
        RECT 0.833000 0.202000 0.923000 0.283000 ;
        RECT 0.451000 0.223000 0.541000 0.304000 ;
        RECT 0.048000 0.195000 0.138000 0.276000 ;
        RECT 0.451000 0.221000 0.526000 0.304000 ;
        RECT 1.214000 0.154000 1.275000 0.256000 ;
        RECT 0.862000 0.154000 0.923000 0.283000 ;
        RECT 0.833000 0.202000 0.894000 0.405000 ;
        RECT 0.480000 0.223000 0.541000 0.405000 ;
        RECT 0.480000 0.350000 0.894000 0.405000 ;
        RECT 0.048000 0.221000 0.526000 0.276000 ;
        RECT 0.862000 0.154000 1.275000 0.208000 ;
        RECT 0.048000 0.223000 0.541000 0.276000 ;
        RECT 0.480000 0.221000 0.526000 0.405000 ;
        RECT 0.862000 0.154000 0.894000 0.405000 ;
    END
END OAI21X2

MACRO OAI211X2
    CLASS CORE ;
    FOREIGN OAI211X2 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 1.800000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.123000 0.426000 0.215000 0.514000 ;
        RECT 0.668000 0.605000 0.761000 0.686000 ;
        RECT 0.123000 0.433000 0.239000 0.514000 ;
        RECT 0.121000 0.439000 0.239000 0.514000 ;
        RECT 0.668000 0.460000 0.731000 0.686000 ;
        RECT 0.059000 0.439000 0.239000 0.494000 ;
        RECT 0.121000 0.460000 0.731000 0.514000 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.333000 0.614000 0.502000 0.707000 ;
        RECT 0.333000 0.614000 0.578000 0.695000 ;
        RECT 0.419000 0.614000 0.487000 0.761000 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.140000 0.426000 1.364000 0.507000 ;
        RECT 1.140000 0.439000 1.381000 0.494000 ;
        END
    END B0
    PIN C0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.475000 0.419000 1.568000 0.500000 ;
        RECT 1.475000 0.419000 1.538000 0.627000 ;
        RECT 0.950000 0.460000 1.013000 0.627000 ;
        RECT 0.950000 0.573000 1.538000 0.627000 ;
        END
    END C0
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 1.800000 1.280000 ;
        RECT 0.976000 1.078000 1.069000 1.280000 ;
        RECT 0.409000 1.078000 0.502000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 1.800000 0.080000 ;
        RECT 0.660000 -0.080000 0.753000 0.280000 ;
        RECT 0.256000 -0.080000 0.349000 0.122000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.769000 0.865000 0.862000 0.952000 ;
        RECT 1.205000 0.283000 1.298000 0.364000 ;
        RECT 1.184000 0.865000 1.320000 0.946000 ;
        RECT 0.049000 0.865000 0.142000 0.946000 ;
        RECT 1.631000 0.310000 1.694000 0.755000 ;
        RECT 1.478000 0.706000 1.541000 0.920000 ;
        RECT 1.499000 0.700000 1.561000 0.761000 ;
        RECT 1.205000 0.306000 1.319000 0.364000 ;
        RECT 1.499000 0.700000 1.694000 0.755000 ;
        RECT 1.478000 0.706000 1.561000 0.761000 ;
        RECT 0.049000 0.865000 1.541000 0.920000 ;
        RECT 1.205000 0.310000 1.694000 0.364000 ;
        RECT 1.499000 0.700000 1.541000 0.920000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 1.555000 0.171000 1.647000 0.252000 ;
        RECT 0.856000 0.202000 0.949000 0.283000 ;
        RECT 0.464000 0.223000 0.556000 0.304000 ;
        RECT 0.049000 0.195000 0.142000 0.276000 ;
        RECT 0.464000 0.221000 0.541000 0.304000 ;
        RECT 0.886000 0.174000 0.949000 0.283000 ;
        RECT 0.856000 0.202000 0.919000 0.405000 ;
        RECT 0.494000 0.223000 0.556000 0.405000 ;
        RECT 0.886000 0.174000 1.647000 0.229000 ;
        RECT 0.494000 0.350000 0.919000 0.405000 ;
        RECT 0.049000 0.221000 0.541000 0.276000 ;
        RECT 0.049000 0.223000 0.556000 0.276000 ;
        RECT 0.494000 0.221000 0.541000 0.405000 ;
        RECT 0.886000 0.174000 0.919000 0.405000 ;
    END
END OAI211X2

MACRO NOR4BBX2
    CLASS CORE ;
    FOREIGN NOR4BBX2 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 2.000000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN AN
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.160000 0.380000 0.249000 0.500000 ;
        RECT 0.160000 0.433000 0.348000 0.500000 ;
        END
    END AN
    PIN BN
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.556000 0.277000 1.780000 0.396000 ;
        END
    END BN
    PIN C
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.501000 0.457000 0.595000 0.538000 ;
        RECT 0.517000 0.457000 0.595000 0.758000 ;
        RECT 1.315000 0.570000 1.379000 0.758000 ;
        RECT 1.332000 0.704000 1.395000 0.761000 ;
        RECT 1.315000 0.570000 1.416000 0.625000 ;
        RECT 0.517000 0.704000 1.395000 0.758000 ;
        RECT 1.332000 0.570000 1.379000 0.761000 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.315000 0.557000 0.379000 0.876000 ;
        RECT 1.500000 0.570000 1.563000 0.876000 ;
        RECT 0.423000 0.821000 0.486000 0.894000 ;
        RECT 1.500000 0.570000 1.602000 0.625000 ;
        RECT 0.315000 0.821000 1.563000 0.876000 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 2.000000 1.280000 ;
        RECT 0.204000 1.078000 0.298000 1.280000 ;
        RECT 1.590000 1.078000 1.683000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 2.000000 0.080000 ;
        RECT 1.074000 -0.080000 1.168000 0.122000 ;
        RECT 0.248000 -0.080000 0.342000 0.198000 ;
        RECT 0.656000 -0.080000 0.749000 0.122000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.857000 0.894000 1.964000 0.986000 ;
        RECT 0.917000 0.931000 1.032000 1.012000 ;
        RECT 0.865000 0.165000 0.959000 0.246000 ;
        RECT 0.446000 0.165000 0.540000 0.246000 ;
        RECT 1.231000 0.150000 1.295000 0.246000 ;
        RECT 0.968000 0.931000 1.032000 1.027000 ;
        RECT 1.901000 0.150000 1.964000 0.986000 ;
        RECT 1.231000 0.150000 1.964000 0.205000 ;
        RECT 0.917000 0.931000 1.964000 0.986000 ;
        RECT 0.446000 0.192000 1.295000 0.246000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 0.033000 0.683000 0.143000 0.876000 ;
        RECT 0.033000 0.217000 0.143000 0.324000 ;
        RECT 1.138000 0.457000 1.231000 0.538000 ;
        RECT 0.919000 0.457000 1.012000 0.538000 ;
        RECT 0.697000 0.457000 0.791000 0.538000 ;
        RECT 0.727000 0.457000 0.791000 0.649000 ;
        RECT 0.318000 0.269000 0.382000 0.379000 ;
        RECT 1.774000 0.457000 1.837000 0.764000 ;
        RECT 1.358000 0.262000 1.421000 0.512000 ;
        RECT 1.138000 0.457000 1.201000 0.649000 ;
        RECT 0.919000 0.324000 0.982000 0.538000 ;
        RECT 0.033000 0.217000 0.096000 0.876000 ;
        RECT 1.358000 0.262000 1.493000 0.317000 ;
        RECT 1.138000 0.457000 1.837000 0.512000 ;
        RECT 0.727000 0.594000 1.201000 0.649000 ;
        RECT 0.318000 0.324000 0.982000 0.379000 ;
        RECT 0.143000 0.269000 0.382000 0.324000 ;
    END
END NOR4BBX2

MACRO NOR4BX2
    CLASS CORE ;
    FOREIGN NOR4BX2 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 1.800000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN AN
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.160000 0.433000 0.322000 0.513000 ;
        RECT 0.160000 0.395000 0.222000 0.513000 ;
        END
    END AN
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.139000 0.452000 1.276000 0.627000 ;
        RECT 0.747000 0.452000 0.840000 0.533000 ;
        RECT 0.747000 0.452000 1.276000 0.507000 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.400000 0.396000 1.561000 0.500000 ;
        RECT 0.578000 0.343000 0.682000 0.439000 ;
        RECT 1.400000 0.343000 1.480000 0.500000 ;
        RECT 0.578000 0.343000 0.641000 0.533000 ;
        RECT 0.578000 0.343000 1.480000 0.398000 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.297000 0.569000 0.390000 0.761000 ;
        RECT 1.519000 0.557000 1.612000 0.638000 ;
        RECT 1.518000 0.570000 1.612000 0.638000 ;
        RECT 1.518000 0.570000 1.580000 0.761000 ;
        RECT 1.519000 0.557000 1.580000 0.761000 ;
        RECT 0.297000 0.700000 0.419000 0.761000 ;
        RECT 0.297000 0.706000 1.580000 0.761000 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 1.800000 1.280000 ;
        RECT 1.631000 1.078000 1.724000 1.280000 ;
        RECT 0.235000 1.078000 0.327000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 1.800000 0.080000 ;
        RECT 0.649000 -0.080000 0.742000 0.122000 ;
        RECT 0.245000 -0.080000 0.338000 0.198000 ;
        RECT 1.064000 -0.080000 1.156000 0.122000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.965000 0.826000 1.058000 0.907000 ;
        RECT 0.856000 0.179000 0.949000 0.260000 ;
        RECT 1.658000 0.192000 1.737000 0.306000 ;
        RECT 0.965000 0.833000 1.140000 0.900000 ;
        RECT 1.675000 0.192000 1.737000 0.894000 ;
        RECT 0.965000 0.839000 1.737000 0.894000 ;
        RECT 0.442000 0.192000 1.737000 0.246000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 0.034000 0.683000 0.142000 0.876000 ;
        RECT 0.034000 0.217000 0.142000 0.323000 ;
        RECT 0.926000 0.570000 1.023000 0.643000 ;
        RECT 0.296000 0.268000 0.359000 0.356000 ;
        RECT 0.034000 0.217000 0.097000 0.876000 ;
        RECT 0.453000 0.301000 0.515000 0.643000 ;
        RECT 0.453000 0.588000 1.023000 0.643000 ;
        RECT 0.296000 0.301000 0.515000 0.356000 ;
        RECT 0.142000 0.268000 0.359000 0.323000 ;
    END
END NOR4BX2

MACRO NOR4X4
    CLASS CORE ;
    FOREIGN NOR4X4 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 3.000000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.691000 0.573000 0.858000 0.679000 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.864000 0.433000 1.999000 0.538000 ;
        RECT 0.512000 0.392000 0.648000 0.494000 ;
        RECT 1.000000 0.392000 1.091000 0.637000 ;
        RECT 0.512000 0.392000 0.603000 0.538000 ;
        RECT 2.352000 0.457000 2.443000 0.538000 ;
        RECT 1.864000 0.392000 1.925000 0.538000 ;
        RECT 1.864000 0.483000 2.443000 0.538000 ;
        RECT 0.512000 0.392000 1.925000 0.446000 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 2.531000 0.476000 2.622000 0.573000 ;
        RECT 1.178000 0.700000 1.262000 0.789000 ;
        RECT 0.362000 0.706000 0.472000 0.789000 ;
        RECT 1.626000 0.502000 1.754000 0.583000 ;
        RECT 1.201000 0.502000 1.291000 0.583000 ;
        RECT 0.333000 0.556000 0.424000 0.637000 ;
        RECT 0.362000 0.556000 0.424000 0.789000 ;
        RECT 2.531000 0.476000 2.592000 0.648000 ;
        RECT 1.693000 0.502000 1.754000 0.648000 ;
        RECT 1.201000 0.502000 1.262000 0.789000 ;
        RECT 1.693000 0.593000 2.592000 0.648000 ;
        RECT 1.201000 0.502000 1.754000 0.557000 ;
        RECT 0.362000 0.735000 1.262000 0.789000 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.425000 0.618000 1.516000 0.758000 ;
        RECT 2.710000 0.429000 2.809000 0.510000 ;
        RECT 0.055000 0.556000 0.237000 0.637000 ;
        RECT 1.425000 0.618000 1.487000 0.899000 ;
        RECT 0.175000 0.556000 0.237000 0.899000 ;
        RECT 2.710000 0.429000 2.771000 0.758000 ;
        RECT 0.175000 0.844000 1.487000 0.899000 ;
        RECT 1.425000 0.704000 2.771000 0.758000 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 3.000000 1.280000 ;
        RECT 1.432000 1.078000 1.523000 1.280000 ;
        RECT 0.048000 1.078000 0.139000 1.280000 ;
        RECT 2.816000 1.078000 2.906000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 3.000000 0.080000 ;
        RECT 2.424000 -0.080000 2.515000 0.212000 ;
        RECT 2.037000 -0.080000 2.128000 0.212000 ;
        RECT 0.834000 -0.080000 0.925000 0.212000 ;
        RECT 0.440000 -0.080000 0.531000 0.211000 ;
        RECT 0.048000 -0.080000 0.139000 0.211000 ;
        RECT 2.816000 -0.080000 2.906000 0.212000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 2.861000 0.567000 2.963000 0.900000 ;
        RECT 2.861000 0.567000 2.943000 0.923000 ;
        RECT 2.619000 0.256000 2.710000 0.337000 ;
        RECT 2.230000 0.256000 2.321000 0.337000 ;
        RECT 2.108000 0.867000 2.199000 0.948000 ;
        RECT 0.755000 0.954000 0.846000 1.035000 ;
        RECT 0.638000 0.256000 0.729000 0.337000 ;
        RECT 0.245000 0.256000 0.336000 0.337000 ;
        RECT 2.881000 0.282000 2.943000 0.923000 ;
        RECT 2.108000 0.867000 2.170000 1.008000 ;
        RECT 2.108000 0.868000 2.943000 0.923000 ;
        RECT 0.245000 0.282000 2.943000 0.337000 ;
        RECT 0.755000 0.954000 2.170000 1.008000 ;
        END
    END Y
END NOR4X4

MACRO NOR4X2
    CLASS CORE ;
    FOREIGN NOR4X2 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 1.600000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.710000 0.555000 0.878000 0.636000 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.517000 0.439000 0.607000 0.538000 ;
        RECT 1.007000 0.556000 1.099000 0.637000 ;
        RECT 0.516000 0.457000 0.607000 0.538000 ;
        RECT 1.007000 0.444000 1.069000 0.637000 ;
        RECT 0.517000 0.439000 0.653000 0.499000 ;
        RECT 0.517000 0.444000 1.069000 0.499000 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.365000 0.706000 0.475000 0.789000 ;
        RECT 1.145000 0.396000 1.236000 0.477000 ;
        RECT 0.335000 0.556000 0.427000 0.637000 ;
        RECT 1.174000 0.396000 1.236000 0.789000 ;
        RECT 0.365000 0.556000 0.427000 0.789000 ;
        RECT 0.365000 0.735000 1.236000 0.789000 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.325000 0.556000 1.417000 0.637000 ;
        RECT 0.055000 0.556000 0.238000 0.637000 ;
        RECT 1.325000 0.556000 1.387000 0.899000 ;
        RECT 0.176000 0.556000 0.238000 0.899000 ;
        RECT 0.176000 0.844000 1.387000 0.899000 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 1.600000 1.280000 ;
        RECT 1.442000 1.078000 1.534000 1.280000 ;
        RECT 0.048000 1.078000 0.140000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 1.600000 0.080000 ;
        RECT 0.501000 -0.080000 0.593000 0.122000 ;
        RECT 0.048000 -0.080000 0.140000 0.225000 ;
        RECT 0.927000 -0.080000 1.018000 0.122000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.460000 0.894000 1.542000 1.008000 ;
        RECT 0.761000 0.954000 0.853000 1.035000 ;
        RECT 0.722000 0.261000 0.813000 0.342000 ;
        RECT 0.246000 0.261000 0.338000 0.342000 ;
        RECT 1.480000 0.287000 1.542000 1.008000 ;
        RECT 0.246000 0.287000 1.542000 0.342000 ;
        RECT 0.761000 0.954000 1.542000 1.008000 ;
        END
    END Y
END NOR4X2

MACRO NOR3BX4
    CLASS CORE ;
    FOREIGN NOR3BX4 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 2.000000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN AN
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.180000 0.438000 0.284000 0.519000 ;
        RECT 0.220000 0.306000 0.284000 0.519000 ;
        RECT 0.220000 0.306000 0.304000 0.361000 ;
        END
    END AN
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.565000 0.411000 0.668000 0.513000 ;
        RECT 0.565000 0.411000 0.658000 0.514000 ;
        RECT 1.034000 0.520000 1.128000 0.606000 ;
        RECT 1.032000 0.411000 1.098000 0.500000 ;
        RECT 1.034000 0.411000 1.098000 0.606000 ;
        RECT 1.561000 0.523000 1.624000 0.606000 ;
        RECT 1.034000 0.551000 1.624000 0.606000 ;
        RECT 0.565000 0.411000 1.098000 0.465000 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.231000 0.414000 1.455000 0.495000 ;
        RECT 0.366000 0.536000 0.486000 0.617000 ;
        RECT 1.231000 0.301000 1.295000 0.495000 ;
        RECT 0.423000 0.301000 0.486000 0.627000 ;
        RECT 0.423000 0.301000 1.295000 0.356000 ;
        END
    END C
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 2.000000 1.280000 ;
        RECT 0.264000 0.866000 0.358000 1.280000 ;
        RECT 1.295000 0.911000 1.388000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 2.000000 0.080000 ;
        RECT 1.128000 -0.080000 1.222000 0.122000 ;
        RECT 0.708000 -0.080000 0.802000 0.122000 ;
        RECT 0.300000 -0.080000 0.394000 0.198000 ;
        RECT 1.536000 -0.080000 1.629000 0.198000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.857000 0.433000 1.961000 0.852000 ;
        RECT 1.807000 0.771000 1.961000 0.852000 ;
        RECT 1.337000 0.165000 1.431000 0.246000 ;
        RECT 0.917000 0.165000 1.011000 0.246000 ;
        RECT 0.782000 0.812000 0.876000 0.893000 ;
        RECT 0.499000 0.165000 0.592000 0.246000 ;
        RECT 0.968000 0.771000 1.052000 0.839000 ;
        RECT 0.968000 0.771000 1.032000 0.867000 ;
        RECT 1.857000 0.268000 1.920000 0.852000 ;
        RECT 1.368000 0.165000 1.431000 0.323000 ;
        RECT 1.368000 0.268000 1.920000 0.323000 ;
        RECT 0.968000 0.771000 1.961000 0.826000 ;
        RECT 0.782000 0.812000 1.032000 0.867000 ;
        RECT 0.499000 0.192000 1.431000 0.246000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 0.780000 0.520000 0.879000 0.756000 ;
        RECT 0.050000 0.701000 0.143000 0.790000 ;
        RECT 0.050000 0.198000 0.157000 0.282000 ;
        RECT 1.687000 0.377000 1.769000 0.715000 ;
        RECT 0.050000 0.198000 0.113000 0.790000 ;
        RECT 1.667000 0.377000 1.769000 0.437000 ;
        RECT 0.050000 0.701000 0.879000 0.756000 ;
        RECT 0.780000 0.661000 1.769000 0.715000 ;
    END
END NOR3BX4

MACRO NOR3BX2
    CLASS CORE ;
    FOREIGN NOR3BX2 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 1.400000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN AN
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.174000 0.376000 0.273000 0.457000 ;
        RECT 0.212000 0.306000 0.273000 0.457000 ;
        RECT 0.212000 0.306000 0.293000 0.361000 ;
        END
    END AN
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.996000 0.555000 1.086000 0.636000 ;
        RECT 0.558000 0.439000 0.643000 0.515000 ;
        RECT 0.996000 0.461000 1.057000 0.636000 ;
        RECT 0.558000 0.439000 0.619000 0.542000 ;
        RECT 0.558000 0.461000 1.057000 0.515000 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.365000 0.536000 0.467000 0.627000 ;
        RECT 1.119000 0.394000 1.209000 0.475000 ;
        RECT 0.335000 0.536000 0.467000 0.617000 ;
        RECT 0.387000 0.494000 0.467000 0.627000 ;
        RECT 1.119000 0.324000 1.180000 0.475000 ;
        RECT 0.406000 0.324000 0.467000 0.627000 ;
        RECT 0.406000 0.324000 1.180000 0.379000 ;
        RECT 0.365000 0.573000 0.468000 0.627000 ;
        END
    END C
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 1.400000 1.280000 ;
        RECT 1.246000 0.932000 1.336000 1.280000 ;
        RECT 0.255000 0.897000 0.345000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 1.400000 0.080000 ;
        RECT 0.681000 -0.080000 0.772000 0.122000 ;
        RECT 0.289000 -0.080000 0.379000 0.198000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.753000 0.806000 0.843000 0.895000 ;
        RECT 0.883000 0.165000 0.973000 0.246000 ;
        RECT 0.480000 0.165000 0.570000 0.246000 ;
        RECT 1.262000 0.761000 1.331000 0.861000 ;
        RECT 1.262000 0.192000 1.331000 0.306000 ;
        RECT 1.270000 0.192000 1.331000 0.861000 ;
        RECT 0.932000 0.806000 0.993000 0.894000 ;
        RECT 0.753000 0.806000 1.331000 0.861000 ;
        RECT 0.480000 0.192000 1.331000 0.246000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 0.048000 0.198000 0.151000 0.282000 ;
        RECT 0.048000 0.670000 0.138000 0.751000 ;
        RECT 0.785000 0.570000 0.846000 0.751000 ;
        RECT 0.048000 0.198000 0.109000 0.751000 ;
        RECT 0.785000 0.570000 0.875000 0.625000 ;
        RECT 0.048000 0.696000 0.846000 0.751000 ;
    END
END NOR3BX2

MACRO NOR3X4
    CLASS CORE ;
    FOREIGN NOR3X4 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 1.800000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.638000 0.379000 0.731000 0.496000 ;
        RECT 1.489000 0.581000 1.582000 0.662000 ;
        RECT 0.599000 0.429000 0.731000 0.494000 ;
        RECT 1.490000 0.379000 1.553000 0.662000 ;
        RECT 0.638000 0.379000 1.553000 0.433000 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.311000 0.507000 0.404000 0.610000 ;
        RECT 0.908000 0.488000 0.971000 0.610000 ;
        RECT 0.311000 0.439000 0.374000 0.610000 ;
        RECT 0.908000 0.488000 1.390000 0.543000 ;
        RECT 0.311000 0.555000 0.971000 0.610000 ;
        RECT 0.239000 0.439000 0.374000 0.494000 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.092000 0.598000 1.189000 0.774000 ;
        RECT 0.056000 0.526000 0.153000 0.627000 ;
        RECT 1.021000 0.700000 1.189000 0.774000 ;
        RECT 0.090000 0.526000 0.153000 0.774000 ;
        RECT 0.090000 0.719000 1.189000 0.774000 ;
        END
    END C
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 1.800000 1.280000 ;
        RECT 1.088000 0.989000 1.181000 1.280000 ;
        RECT 0.049000 0.929000 0.142000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 1.800000 0.080000 ;
        RECT 1.227000 -0.080000 1.320000 0.198000 ;
        RECT 0.442000 -0.080000 0.535000 0.198000 ;
        RECT 0.049000 -0.080000 0.142000 0.211000 ;
        RECT 0.835000 -0.080000 0.927000 0.198000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.658000 0.567000 1.762000 0.900000 ;
        RECT 1.561000 0.810000 1.762000 0.892000 ;
        RECT 1.031000 0.242000 1.124000 0.323000 ;
        RECT 0.638000 0.242000 0.731000 0.323000 ;
        RECT 0.573000 0.837000 0.665000 0.918000 ;
        RECT 0.245000 0.242000 0.338000 0.323000 ;
        RECT 1.658000 0.268000 1.721000 0.900000 ;
        RECT 0.573000 0.837000 1.762000 0.892000 ;
        RECT 0.245000 0.268000 1.721000 0.323000 ;
        END
    END Y
END NOR3X4

MACRO NOR3X2
    CLASS CORE ;
    FOREIGN NOR3X2 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 1.300000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.498000 0.439000 0.682000 0.525000 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.321000 0.445000 0.415000 0.539000 ;
        RECT 0.847000 0.377000 0.943000 0.458000 ;
        RECT 0.321000 0.458000 0.416000 0.539000 ;
        RECT 0.848000 0.377000 0.913000 0.635000 ;
        RECT 0.352000 0.458000 0.416000 0.635000 ;
        RECT 0.352000 0.445000 0.415000 0.635000 ;
        RECT 0.246000 0.439000 0.311000 0.500000 ;
        RECT 0.352000 0.580000 0.913000 0.635000 ;
        RECT 0.246000 0.445000 0.415000 0.500000 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.118000 0.573000 0.214000 0.707000 ;
        RECT 1.007000 0.537000 1.088000 0.744000 ;
        RECT 0.149000 0.573000 0.214000 0.744000 ;
        RECT 0.149000 0.689000 1.088000 0.744000 ;
        RECT 0.058000 0.573000 0.214000 0.627000 ;
        END
    END C
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 1.300000 1.280000 ;
        RECT 1.109000 0.925000 1.204000 1.280000 ;
        RECT 0.051000 0.876000 0.146000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 1.300000 0.080000 ;
        RECT 0.456000 -0.080000 0.552000 0.211000 ;
        RECT 0.051000 -0.080000 0.146000 0.211000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.658000 0.151000 0.754000 0.344000 ;
        RECT 0.253000 0.151000 0.349000 0.344000 ;
        RECT 0.591000 0.800000 0.687000 0.890000 ;
        RECT 1.154000 0.767000 1.240000 0.855000 ;
        RECT 1.175000 0.255000 1.240000 0.855000 ;
        RECT 0.658000 0.255000 1.240000 0.310000 ;
        RECT 0.591000 0.800000 1.240000 0.855000 ;
        RECT 0.253000 0.289000 0.754000 0.344000 ;
        END
    END Y
END NOR3X2

MACRO NOR2BX4
    CLASS CORE ;
    FOREIGN NOR2BX4 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 1.400000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN AN
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.034000 0.436000 0.138000 0.571000 ;
        END
    END AN
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.321000 0.521000 0.411000 0.650000 ;
        RECT 0.936000 0.563000 1.026000 0.650000 ;
        RECT 0.321000 0.565000 0.468000 0.650000 ;
        RECT 0.321000 0.595000 1.026000 0.650000 ;
        END
    END B
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.223000 1.117000 1.013000 1.280000 ;
        RECT 0.000000 1.120000 1.400000 1.280000 ;
        RECT 0.923000 1.078000 1.013000 1.280000 ;
        RECT 0.223000 1.078000 0.313000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 1.400000 0.080000 ;
        RECT 0.681000 -0.080000 0.772000 0.122000 ;
        RECT 1.087000 -0.080000 1.177000 0.122000 ;
        RECT 0.276000 -0.080000 0.366000 0.122000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.262000 0.264000 1.363000 0.786000 ;
        RECT 1.252000 0.693000 1.363000 0.786000 ;
        RECT 0.883000 0.255000 0.973000 0.336000 ;
        RECT 0.573000 0.705000 1.363000 0.786000 ;
        RECT 0.480000 0.255000 0.570000 0.336000 ;
        RECT 0.883000 0.264000 1.363000 0.336000 ;
        RECT 0.480000 0.281000 1.363000 0.336000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 0.578000 0.392000 0.668000 0.538000 ;
        RECT 0.074000 0.281000 0.164000 0.362000 ;
        RECT 0.048000 0.793000 0.138000 0.874000 ;
        RECT 1.139000 0.392000 1.200000 0.546000 ;
        RECT 0.199000 0.307000 0.260000 0.848000 ;
        RECT 0.074000 0.307000 0.260000 0.362000 ;
        RECT 0.048000 0.793000 0.260000 0.848000 ;
        RECT 0.578000 0.392000 1.200000 0.446000 ;
        RECT 0.260000 0.392000 0.578000 0.446000 ;
    END
END NOR2BX4

MACRO NOR2BX2
    CLASS CORE ;
    FOREIGN NOR2BX2 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 1.100000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN AN
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.050000 0.457000 0.144000 0.633000 ;
        END
    END AN
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.406000 0.300000 0.511000 0.473000 ;
        RECT 0.847000 0.418000 0.928000 0.565000 ;
        RECT 0.342000 0.433000 0.436000 0.514000 ;
        RECT 0.357000 0.418000 0.436000 0.514000 ;
        RECT 0.357000 0.418000 0.928000 0.473000 ;
        RECT 0.406000 0.300000 0.436000 0.514000 ;
        END
    END B
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 1.100000 1.280000 ;
        RECT 0.956000 1.078000 1.050000 1.280000 ;
        RECT 0.228000 1.078000 0.322000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 1.100000 0.080000 ;
        RECT 0.956000 -0.080000 1.050000 0.228000 ;
        RECT 0.542000 -0.080000 0.636000 0.122000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.756000 0.282000 0.850000 0.363000 ;
        RECT 0.594000 0.712000 0.689000 0.793000 ;
        RECT 0.997000 0.308000 1.061000 0.767000 ;
        RECT 0.976000 0.706000 1.061000 0.767000 ;
        RECT 0.756000 0.308000 1.061000 0.363000 ;
        RECT 0.594000 0.712000 1.061000 0.767000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 0.622000 0.538000 0.717000 0.626000 ;
        RECT 0.050000 0.748000 0.144000 0.829000 ;
        RECT 0.050000 0.286000 0.144000 0.367000 ;
        RECT 0.208000 0.312000 0.272000 0.802000 ;
        RECT 0.208000 0.571000 0.717000 0.626000 ;
        RECT 0.050000 0.312000 0.272000 0.367000 ;
        RECT 0.050000 0.748000 0.272000 0.802000 ;
    END
END NOR2BX2

MACRO NOR2X4
    CLASS CORE ;
    FOREIGN NOR2X4 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 1.300000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.432000 0.439000 0.523000 0.525000 ;
        RECT 0.990000 0.464000 1.086000 0.545000 ;
        RECT 0.990000 0.394000 1.055000 0.545000 ;
        RECT 0.459000 0.394000 0.523000 0.525000 ;
        RECT 0.459000 0.394000 1.055000 0.449000 ;
        RECT 0.428000 0.470000 0.523000 0.525000 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.763000 0.561000 0.858000 0.642000 ;
        RECT 0.138000 0.492000 0.234000 0.573000 ;
        RECT 0.246000 0.650000 0.311000 0.761000 ;
        RECT 0.169000 0.492000 0.234000 0.707000 ;
        RECT 0.763000 0.561000 0.827000 0.705000 ;
        RECT 0.169000 0.650000 0.311000 0.707000 ;
        RECT 0.169000 0.650000 0.827000 0.705000 ;
        END
    END B
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 1.300000 1.280000 ;
        RECT 0.799000 1.078000 0.895000 1.280000 ;
        RECT 0.056000 1.078000 0.152000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 1.300000 0.080000 ;
        RECT 0.467000 -0.080000 0.563000 0.211000 ;
        RECT 0.884000 -0.080000 0.979000 0.122000 ;
        RECT 0.051000 -0.080000 0.146000 0.298000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.154000 0.433000 1.261000 0.767000 ;
        RECT 1.148000 0.693000 1.244000 0.840000 ;
        RECT 1.154000 0.433000 1.244000 0.840000 ;
        RECT 1.165000 0.265000 1.249000 0.767000 ;
        RECT 0.670000 0.256000 0.765000 0.337000 ;
        RECT 0.265000 0.256000 0.360000 0.337000 ;
        RECT 0.428000 0.760000 1.244000 0.840000 ;
        RECT 1.165000 0.265000 1.244000 0.840000 ;
        RECT 1.148000 0.693000 1.261000 0.767000 ;
        RECT 0.670000 0.265000 1.249000 0.337000 ;
        RECT 0.265000 0.282000 1.249000 0.337000 ;
        END
    END Y
END NOR2X4

MACRO NOR2X2
    CLASS CORE ;
    FOREIGN NOR2X2 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 0.900000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.327000 0.538000 0.502000 0.633000 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.120000 0.418000 0.229000 0.518000 ;
        RECT 0.652000 0.418000 0.742000 0.564000 ;
        RECT 0.059000 0.418000 0.229000 0.494000 ;
        RECT 0.059000 0.418000 0.742000 0.473000 ;
        END
    END B
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 0.900000 1.280000 ;
        RECT 0.758000 1.078000 0.851000 1.280000 ;
        RECT 0.049000 1.078000 0.142000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 0.900000 0.080000 ;
        RECT 0.758000 -0.080000 0.851000 0.228000 ;
        RECT 0.365000 -0.080000 0.458000 0.340000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.562000 0.170000 0.655000 0.363000 ;
        RECT 0.404000 0.712000 0.496000 0.793000 ;
        RECT 0.805000 0.308000 0.867000 0.761000 ;
        RECT 0.779000 0.706000 0.862000 0.767000 ;
        RECT 0.805000 0.308000 0.862000 0.767000 ;
        RECT 0.779000 0.706000 0.867000 0.761000 ;
        RECT 0.562000 0.308000 0.867000 0.363000 ;
        RECT 0.404000 0.712000 0.862000 0.767000 ;
        END
    END Y
END NOR2X2

MACRO NAND4BBX2
    CLASS CORE ;
    FOREIGN NAND4BBX2 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 2.000000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN AN
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.043000 0.433000 0.147000 0.574000 ;
        END
    END AN
    PIN BN
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.657000 0.498000 1.780000 0.633000 ;
        END
    END BN
    PIN C
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.287000 0.519000 1.380000 0.627000 ;
        RECT 0.522000 0.519000 0.634000 0.600000 ;
        RECT 0.570000 0.519000 0.634000 0.706000 ;
        RECT 1.287000 0.519000 1.350000 0.706000 ;
        RECT 0.570000 0.651000 1.350000 0.706000 ;
        RECT 1.287000 0.573000 1.395000 0.627000 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.365000 0.706000 0.486000 0.815000 ;
        RECT 1.371000 0.761000 1.464000 0.842000 ;
        RECT 0.340000 0.519000 0.428000 0.600000 ;
        RECT 0.365000 0.519000 0.428000 0.815000 ;
        RECT 0.365000 0.761000 1.464000 0.815000 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 2.000000 1.280000 ;
        RECT 1.737000 1.078000 1.882000 1.280000 ;
        RECT 1.017000 1.078000 1.140000 1.280000 ;
        RECT 0.639000 1.078000 0.733000 1.280000 ;
        RECT 0.248000 1.078000 0.342000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.092000 -0.080000 0.318000 0.122000 ;
        RECT 0.000000 -0.080000 2.000000 0.080000 ;
        RECT 1.569000 -0.080000 1.663000 0.122000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.897000 0.150000 0.990000 0.343000 ;
        RECT 0.972000 0.870000 1.055000 0.973000 ;
        RECT 1.879000 0.573000 1.961000 0.973000 ;
        RECT 1.857000 0.893000 1.961000 0.973000 ;
        RECT 1.884000 0.195000 1.961000 0.973000 ;
        RECT 0.972000 0.901000 1.961000 0.973000 ;
        RECT 0.444000 0.870000 1.055000 0.942000 ;
        RECT 1.868000 0.573000 1.961000 0.644000 ;
        RECT 0.897000 0.195000 1.961000 0.262000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 0.050000 0.675000 0.143000 0.868000 ;
        RECT 0.895000 0.400000 0.999000 0.487000 ;
        RECT 1.096000 0.514000 1.200000 0.596000 ;
        RECT 1.528000 0.761000 1.621000 0.842000 ;
        RECT 0.705000 0.515000 0.809000 0.596000 ;
        RECT 0.050000 0.276000 0.143000 0.357000 ;
        RECT 1.528000 0.330000 1.821000 0.398000 ;
        RECT 1.136000 0.401000 1.200000 0.596000 ;
        RECT 1.758000 0.317000 1.821000 0.398000 ;
        RECT 1.528000 0.330000 1.591000 0.842000 ;
        RECT 0.211000 0.302000 0.274000 0.730000 ;
        RECT 1.136000 0.401000 1.591000 0.456000 ;
        RECT 0.705000 0.400000 0.999000 0.455000 ;
        RECT 0.274000 0.400000 0.895000 0.455000 ;
        RECT 0.211000 0.400000 0.809000 0.455000 ;
        RECT 0.050000 0.675000 0.274000 0.730000 ;
        RECT 0.050000 0.302000 0.274000 0.357000 ;
        RECT 0.705000 0.542000 1.200000 0.596000 ;
    END
END NAND4BBX2

MACRO NAND4BX4
    CLASS CORE ;
    FOREIGN NAND4BX4 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 3.200000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN AN
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.042000 0.433000 0.144000 0.574000 ;
        END
    END AN
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 2.349000 0.433000 2.451000 0.596000 ;
        RECT 2.003000 0.510000 2.104000 0.596000 ;
        RECT 1.121000 0.510000 1.222000 0.596000 ;
        RECT 2.349000 0.515000 2.465000 0.596000 ;
        RECT 0.723000 0.515000 0.824000 0.596000 ;
        RECT 2.003000 0.542000 2.465000 0.596000 ;
        RECT 1.121000 0.510000 2.104000 0.564000 ;
        RECT 0.723000 0.542000 1.222000 0.596000 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 2.591000 0.519000 2.683000 0.600000 ;
        RECT 1.825000 0.625000 1.916000 0.706000 ;
        RECT 1.309000 0.625000 1.401000 0.706000 ;
        RECT 0.544000 0.519000 0.653000 0.600000 ;
        RECT 2.591000 0.519000 2.668000 0.633000 ;
        RECT 2.527000 0.579000 2.589000 0.706000 ;
        RECT 0.591000 0.519000 0.653000 0.706000 ;
        RECT 2.547000 0.573000 2.668000 0.633000 ;
        RECT 1.825000 0.651000 2.589000 0.706000 ;
        RECT 1.309000 0.625000 1.916000 0.680000 ;
        RECT 0.591000 0.651000 1.401000 0.706000 ;
        RECT 2.527000 0.579000 2.668000 0.633000 ;
        RECT 2.547000 0.573000 2.589000 0.706000 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 2.769000 0.426000 2.859000 0.507000 ;
        RECT 0.361000 0.519000 0.453000 0.600000 ;
        RECT 1.568000 0.735000 1.659000 0.815000 ;
        RECT 2.753000 0.439000 2.859000 0.507000 ;
        RECT 2.753000 0.439000 2.815000 0.815000 ;
        RECT 0.413000 0.706000 0.475000 0.815000 ;
        RECT 0.391000 0.519000 0.453000 0.761000 ;
        RECT 0.391000 0.706000 0.475000 0.761000 ;
        RECT 0.413000 0.761000 2.815000 0.815000 ;
        RECT 2.769000 0.426000 2.815000 0.815000 ;
        RECT 0.413000 0.519000 0.453000 0.815000 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 3.200000 1.280000 ;
        RECT 2.078000 1.078000 2.199000 1.280000 ;
        RECT 1.028000 1.078000 1.149000 1.280000 ;
        RECT 2.859000 1.078000 2.951000 1.280000 ;
        RECT 0.276000 1.078000 0.368000 1.280000 ;
        RECT 2.477000 1.078000 2.568000 1.280000 ;
        RECT 0.659000 1.078000 0.750000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 3.200000 0.080000 ;
        RECT 2.882000 -0.080000 2.974000 0.122000 ;
        RECT 0.253000 -0.080000 0.345000 0.122000 ;
        RECT 1.568000 -0.080000 1.659000 0.122000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 2.882000 0.567000 2.985000 0.900000 ;
        RECT 2.882000 0.567000 2.974000 0.942000 ;
        RECT 0.910000 0.150000 1.002000 0.343000 ;
        RECT 2.225000 0.150000 2.316000 0.343000 ;
        RECT 2.294000 0.870000 2.974000 0.942000 ;
        RECT 0.910000 0.207000 2.316000 0.274000 ;
        RECT 0.467000 0.870000 2.974000 0.937000 ;
        RECT 2.921000 0.288000 2.983000 0.900000 ;
        RECT 2.225000 0.288000 2.983000 0.343000 ;
        RECT 2.921000 0.288000 2.974000 0.942000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 2.180000 0.400000 2.281000 0.487000 ;
        RECT 0.909000 0.400000 1.010000 0.487000 ;
        RECT 0.048000 0.801000 0.140000 0.882000 ;
        RECT 0.048000 0.276000 0.140000 0.357000 ;
        RECT 0.210000 0.302000 0.272000 0.856000 ;
        RECT 0.909000 0.400000 2.281000 0.455000 ;
        RECT 0.272000 0.400000 0.909000 0.455000 ;
        RECT 0.048000 0.801000 0.272000 0.856000 ;
        RECT 0.048000 0.302000 0.272000 0.357000 ;
    END
END NAND4BX4

MACRO NAND4BX2
    CLASS CORE ;
    FOREIGN NAND4BX2 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 1.800000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN AN
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.042000 0.433000 0.146000 0.574000 ;
        END
    END AN
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.085000 0.514000 1.188000 0.596000 ;
        RECT 0.698000 0.515000 0.800000 0.596000 ;
        RECT 1.118000 0.433000 1.188000 0.596000 ;
        RECT 1.118000 0.439000 1.201000 0.494000 ;
        RECT 0.698000 0.542000 1.188000 0.596000 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.285000 0.519000 1.377000 0.627000 ;
        RECT 0.521000 0.519000 0.627000 0.600000 ;
        RECT 1.285000 0.519000 1.347000 0.706000 ;
        RECT 0.565000 0.519000 0.627000 0.706000 ;
        RECT 0.565000 0.651000 1.347000 0.706000 ;
        RECT 1.285000 0.573000 1.381000 0.627000 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.357000 0.761000 1.450000 0.842000 ;
        RECT 0.340000 0.519000 0.424000 0.600000 ;
        RECT 0.361000 0.519000 0.424000 0.761000 ;
        RECT 0.419000 0.706000 0.481000 0.815000 ;
        RECT 0.361000 0.706000 0.481000 0.761000 ;
        RECT 0.419000 0.761000 1.450000 0.815000 ;
        RECT 0.419000 0.519000 0.424000 0.815000 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 1.800000 1.280000 ;
        RECT 1.006000 1.078000 1.129000 1.280000 ;
        RECT 0.245000 1.078000 0.338000 1.280000 ;
        RECT 0.633000 1.078000 0.725000 1.280000 ;
        RECT 0.260000 1.065000 0.323000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 1.800000 0.080000 ;
        RECT 1.560000 -0.080000 1.653000 0.122000 ;
        RECT 0.229000 -0.080000 0.322000 0.122000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.895000 0.150000 0.987000 0.343000 ;
        RECT 1.658000 0.195000 1.741000 0.306000 ;
        RECT 1.658000 0.564000 1.740000 0.973000 ;
        RECT 0.963000 0.870000 1.045000 0.973000 ;
        RECT 1.665000 0.195000 1.741000 0.633000 ;
        RECT 1.665000 0.195000 1.740000 0.973000 ;
        RECT 0.963000 0.901000 1.740000 0.973000 ;
        RECT 0.439000 0.870000 1.045000 0.942000 ;
        RECT 1.658000 0.564000 1.741000 0.633000 ;
        RECT 0.895000 0.195000 1.741000 0.262000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 0.886000 0.400000 0.989000 0.487000 ;
        RECT 0.049000 0.731000 0.142000 0.812000 ;
        RECT 0.049000 0.276000 0.142000 0.357000 ;
        RECT 0.211000 0.302000 0.274000 0.799000 ;
        RECT 0.274000 0.400000 0.886000 0.455000 ;
        RECT 0.049000 0.744000 0.274000 0.799000 ;
        RECT 0.049000 0.302000 0.274000 0.357000 ;
    END
END NAND4BX2

MACRO NAND4X4
    CLASS CORE ;
    FOREIGN NAND4X4 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 3.000000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.988000 0.400000 2.088000 0.487000 ;
        RECT 0.726000 0.400000 0.826000 0.487000 ;
        RECT 0.430000 0.306000 0.492000 0.455000 ;
        RECT 0.430000 0.400000 2.088000 0.455000 ;
        RECT 0.410000 0.306000 0.492000 0.361000 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 2.155000 0.433000 2.257000 0.596000 ;
        RECT 1.811000 0.510000 1.912000 0.596000 ;
        RECT 0.936000 0.510000 1.036000 0.596000 ;
        RECT 2.155000 0.515000 2.270000 0.596000 ;
        RECT 0.541000 0.515000 0.642000 0.596000 ;
        RECT 1.811000 0.542000 2.270000 0.596000 ;
        RECT 0.936000 0.510000 1.912000 0.564000 ;
        RECT 0.541000 0.542000 1.036000 0.596000 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 2.396000 0.519000 2.487000 0.600000 ;
        RECT 1.635000 0.625000 1.726000 0.706000 ;
        RECT 1.123000 0.625000 1.214000 0.706000 ;
        RECT 0.364000 0.519000 0.472000 0.600000 ;
        RECT 2.396000 0.519000 2.472000 0.633000 ;
        RECT 0.410000 0.519000 0.472000 0.706000 ;
        RECT 2.332000 0.579000 2.393000 0.706000 ;
        RECT 2.352000 0.573000 2.472000 0.633000 ;
        RECT 1.635000 0.651000 2.393000 0.706000 ;
        RECT 1.123000 0.625000 1.726000 0.680000 ;
        RECT 0.410000 0.651000 1.214000 0.706000 ;
        RECT 2.332000 0.579000 2.472000 0.633000 ;
        RECT 2.352000 0.573000 2.393000 0.706000 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 2.572000 0.426000 2.662000 0.507000 ;
        RECT 0.182000 0.519000 0.273000 0.600000 ;
        RECT 1.380000 0.735000 1.471000 0.815000 ;
        RECT 2.556000 0.439000 2.662000 0.507000 ;
        RECT 2.556000 0.439000 2.618000 0.815000 ;
        RECT 0.211000 0.519000 0.273000 0.761000 ;
        RECT 0.234000 0.706000 0.295000 0.815000 ;
        RECT 0.211000 0.706000 0.295000 0.761000 ;
        RECT 0.234000 0.761000 2.618000 0.815000 ;
        RECT 2.572000 0.426000 2.618000 0.815000 ;
        RECT 0.234000 0.519000 0.273000 0.815000 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 3.000000 1.280000 ;
        RECT 1.886000 1.078000 2.007000 1.280000 ;
        RECT 0.844000 1.078000 0.964000 1.280000 ;
        RECT 2.662000 1.078000 2.753000 1.280000 ;
        RECT 2.282000 1.078000 2.373000 1.280000 ;
        RECT 0.477000 1.078000 0.568000 1.280000 ;
        RECT 0.098000 1.078000 0.189000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 3.000000 0.080000 ;
        RECT 2.684000 -0.080000 2.775000 0.122000 ;
        RECT 1.380000 -0.080000 1.471000 0.122000 ;
        RECT 0.075000 -0.080000 0.166000 0.122000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 2.684000 0.192000 2.803000 0.307000 ;
        RECT 2.032000 0.150000 2.176000 0.263000 ;
        RECT 2.684000 0.567000 2.786000 0.900000 ;
        RECT 2.684000 0.567000 2.775000 0.942000 ;
        RECT 2.032000 0.150000 2.123000 0.343000 ;
        RECT 0.727000 0.150000 0.818000 0.343000 ;
        RECT 2.723000 0.192000 2.803000 0.639000 ;
        RECT 2.684000 0.567000 2.803000 0.639000 ;
        RECT 2.100000 0.870000 2.775000 0.942000 ;
        RECT 2.032000 0.192000 2.803000 0.263000 ;
        RECT 0.727000 0.207000 2.123000 0.274000 ;
        RECT 0.287000 0.870000 2.775000 0.937000 ;
        RECT 2.723000 0.192000 2.786000 0.900000 ;
        RECT 0.727000 0.207000 2.803000 0.263000 ;
        RECT 2.723000 0.192000 2.775000 0.942000 ;
        END
    END Y
END NAND4X4

MACRO NAND4X2
    CLASS CORE ;
    FOREIGN NAND4X2 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 1.600000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.698000 0.401000 0.799000 0.487000 ;
        RECT 0.434000 0.306000 0.496000 0.456000 ;
        RECT 0.434000 0.401000 0.799000 0.456000 ;
        RECT 0.413000 0.306000 0.496000 0.361000 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.916000 0.439000 1.017000 0.596000 ;
        RECT 0.512000 0.515000 0.613000 0.596000 ;
        RECT 0.512000 0.542000 1.017000 0.596000 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.102000 0.519000 1.187000 0.627000 ;
        RECT 1.102000 0.519000 1.193000 0.600000 ;
        RECT 0.333000 0.519000 0.442000 0.600000 ;
        RECT 1.102000 0.519000 1.164000 0.706000 ;
        RECT 0.380000 0.519000 0.442000 0.706000 ;
        RECT 0.380000 0.651000 1.164000 0.706000 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.162000 0.761000 1.254000 0.842000 ;
        RECT 0.149000 0.519000 0.241000 0.600000 ;
        RECT 0.236000 0.706000 0.298000 0.815000 ;
        RECT 0.179000 0.519000 0.241000 0.761000 ;
        RECT 0.179000 0.706000 0.298000 0.761000 ;
        RECT 0.236000 0.761000 1.254000 0.815000 ;
        RECT 0.236000 0.519000 0.241000 0.815000 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 1.600000 1.280000 ;
        RECT 0.816000 1.078000 0.937000 1.280000 ;
        RECT 0.447000 1.078000 0.539000 1.280000 ;
        RECT 0.065000 1.078000 0.156000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 1.600000 0.080000 ;
        RECT 1.363000 -0.080000 1.455000 0.122000 ;
        RECT 0.048000 -0.080000 0.140000 0.122000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.706000 0.150000 0.797000 0.343000 ;
        RECT 1.460000 0.195000 1.542000 0.306000 ;
        RECT 1.460000 0.564000 1.541000 0.973000 ;
        RECT 0.773000 0.870000 0.854000 0.973000 ;
        RECT 1.467000 0.195000 1.542000 0.633000 ;
        RECT 1.467000 0.195000 1.541000 0.973000 ;
        RECT 0.773000 0.901000 1.541000 0.973000 ;
        RECT 0.256000 0.870000 0.854000 0.942000 ;
        RECT 1.460000 0.564000 1.542000 0.633000 ;
        RECT 0.706000 0.195000 1.542000 0.262000 ;
        END
    END Y
END NAND4X2

MACRO NAND3BX4
    CLASS CORE ;
    FOREIGN NAND3BX4 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 2.000000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN AN
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.047000 0.411000 0.140000 0.563000 ;
        END
    END AN
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.039000 0.507000 1.234000 0.633000 ;
        RECT 1.489000 0.507000 1.583000 0.607000 ;
        RECT 1.039000 0.494000 1.132000 0.633000 ;
        RECT 0.567000 0.577000 0.661000 0.658000 ;
        RECT 1.032000 0.567000 1.234000 0.633000 ;
        RECT 1.039000 0.507000 1.583000 0.562000 ;
        RECT 0.567000 0.579000 1.234000 0.633000 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.234000 0.915000 1.328000 0.996000 ;
        RECT 0.333000 0.439000 0.397000 0.983000 ;
        RECT 0.333000 0.439000 0.486000 0.500000 ;
        RECT 0.333000 0.929000 1.328000 0.983000 ;
        END
    END C
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 2.000000 1.280000 ;
        RECT 1.434000 0.905000 1.528000 1.280000 ;
        RECT 1.070000 1.078000 1.164000 1.280000 ;
        RECT 0.687000 1.078000 0.781000 1.280000 ;
        RECT 0.269000 1.078000 0.362000 1.280000 ;
        RECT 1.843000 0.905000 1.906000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 2.000000 0.080000 ;
        RECT 1.311000 -0.080000 1.405000 0.122000 ;
        RECT 0.264000 -0.080000 0.358000 0.122000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.577000 0.688000 1.723000 0.810000 ;
        RECT 1.577000 0.700000 1.780000 0.810000 ;
        RECT 1.675000 0.700000 1.780000 1.033000 ;
        RECT 1.846000 0.199000 1.950000 0.307000 ;
        RECT 0.788000 0.167000 0.882000 0.254000 ;
        RECT 0.883000 0.742000 0.977000 0.823000 ;
        RECT 0.492000 0.742000 0.585000 0.823000 ;
        RECT 0.850000 0.742000 0.977000 0.810000 ;
        RECT 1.887000 0.199000 1.950000 0.755000 ;
        RECT 1.577000 0.700000 1.950000 0.755000 ;
        RECT 0.788000 0.199000 1.950000 0.254000 ;
        RECT 0.492000 0.755000 1.780000 0.810000 ;
        RECT 1.675000 0.688000 1.723000 1.033000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 0.755000 0.315000 0.848000 0.496000 ;
        RECT 0.050000 0.690000 0.143000 0.771000 ;
        RECT 0.050000 0.224000 0.143000 0.305000 ;
        RECT 1.759000 0.440000 1.822000 0.555000 ;
        RECT 1.712000 0.315000 1.775000 0.495000 ;
        RECT 0.207000 0.250000 0.270000 0.745000 ;
        RECT 1.712000 0.440000 1.822000 0.495000 ;
        RECT 0.755000 0.315000 1.775000 0.370000 ;
        RECT 0.270000 0.315000 0.755000 0.370000 ;
        RECT 0.050000 0.690000 0.270000 0.745000 ;
        RECT 0.050000 0.250000 0.270000 0.305000 ;
        RECT 1.759000 0.315000 1.775000 0.555000 ;
    END
END NAND3BX4

MACRO NAND3BX2
    CLASS CORE ;
    FOREIGN NAND3BX2 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 1.400000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN AN
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.262000 0.467000 1.363000 0.594000 ;
        RECT 1.267000 0.433000 1.358000 0.594000 ;
        END
    END AN
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.737000 0.433000 0.838000 0.604000 ;
        RECT 0.355000 0.514000 0.445000 0.604000 ;
        RECT 0.737000 0.507000 0.870000 0.588000 ;
        RECT 0.355000 0.549000 0.838000 0.604000 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.082000 0.439000 0.172000 0.573000 ;
        RECT 0.957000 0.462000 1.047000 0.543000 ;
        RECT 0.972000 0.462000 1.033000 0.881000 ;
        RECT 0.111000 0.439000 0.172000 0.881000 ;
        RECT 0.111000 0.826000 1.033000 0.881000 ;
        RECT 0.057000 0.439000 0.172000 0.494000 ;
        END
    END C
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 1.400000 1.280000 ;
        RECT 1.058000 0.952000 1.148000 1.280000 ;
        RECT 0.471000 0.952000 0.561000 1.280000 ;
        RECT 0.102000 0.952000 0.192000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 1.400000 0.080000 ;
        RECT 1.055000 -0.080000 1.161000 0.122000 ;
        RECT 1.055000 -0.080000 1.145000 0.247000 ;
        RECT 0.064000 -0.080000 0.154000 0.247000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.651000 0.689000 0.741000 0.770000 ;
        RECT 0.567000 0.164000 0.658000 0.245000 ;
        RECT 0.282000 0.689000 0.373000 0.770000 ;
        RECT 0.643000 0.689000 0.741000 0.767000 ;
        RECT 0.233000 0.689000 0.407000 0.767000 ;
        RECT 0.233000 0.700000 0.741000 0.767000 ;
        RECT 0.233000 0.177000 0.294000 0.767000 ;
        RECT 0.233000 0.177000 0.658000 0.232000 ;
        RECT 0.282000 0.177000 0.294000 0.770000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 1.262000 0.279000 1.352000 0.379000 ;
        RECT 1.262000 0.702000 1.352000 0.783000 ;
        RECT 0.567000 0.410000 0.658000 0.490000 ;
        RECT 1.140000 0.324000 1.201000 0.757000 ;
        RECT 0.597000 0.324000 0.658000 0.490000 ;
        RECT 1.140000 0.702000 1.352000 0.757000 ;
        RECT 0.597000 0.324000 1.352000 0.379000 ;
    END
END NAND3BX2

MACRO NAND3X4
    CLASS CORE ;
    FOREIGN NAND3X4 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 1.800000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.486000 0.426000 1.579000 0.590000 ;
        RECT 0.584000 0.411000 0.676000 0.492000 ;
        RECT 1.484000 0.426000 1.579000 0.499000 ;
        RECT 1.484000 0.302000 1.546000 0.499000 ;
        RECT 0.614000 0.302000 0.676000 0.492000 ;
        RECT 1.486000 0.302000 1.546000 0.590000 ;
        RECT 0.614000 0.302000 1.546000 0.357000 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.302000 0.494000 1.395000 0.590000 ;
        RECT 0.385000 0.514000 0.477000 0.601000 ;
        RECT 0.835000 0.417000 0.927000 0.498000 ;
        RECT 0.758000 0.418000 0.927000 0.498000 ;
        RECT 1.302000 0.418000 1.365000 0.590000 ;
        RECT 0.758000 0.418000 0.821000 0.601000 ;
        RECT 0.758000 0.418000 1.365000 0.473000 ;
        RECT 0.385000 0.546000 0.821000 0.601000 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.059000 0.439000 0.155000 0.573000 ;
        RECT 1.020000 0.527000 1.113000 0.608000 ;
        RECT 1.035000 0.527000 1.098000 0.880000 ;
        RECT 0.093000 0.439000 0.155000 0.880000 ;
        RECT 0.093000 0.825000 1.098000 0.880000 ;
        END
    END C
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 1.800000 1.280000 ;
        RECT 1.602000 0.952000 1.695000 1.280000 ;
        RECT 1.231000 0.952000 1.324000 1.280000 ;
        RECT 0.863000 0.952000 0.956000 1.280000 ;
        RECT 0.484000 0.952000 0.577000 1.280000 ;
        RECT 0.105000 0.952000 0.198000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 1.800000 0.080000 ;
        RECT 1.102000 -0.080000 1.195000 0.122000 ;
        RECT 0.063000 -0.080000 0.155000 0.247000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.218000 0.167000 0.322000 0.500000 ;
        RECT 1.620000 0.158000 1.713000 0.351000 ;
        RECT 0.224000 0.167000 0.316000 0.770000 ;
        RECT 1.560000 0.158000 1.713000 0.248000 ;
        RECT 1.417000 0.689000 1.510000 0.770000 ;
        RECT 0.224000 0.689000 0.770000 0.770000 ;
        RECT 0.218000 0.167000 0.676000 0.248000 ;
        RECT 1.645000 0.158000 1.707000 0.744000 ;
        RECT 1.417000 0.689000 1.707000 0.744000 ;
        RECT 0.218000 0.193000 1.713000 0.248000 ;
        END
    END Y
END NAND3X4

MACRO NAND3X2
    CLASS CORE ;
    FOREIGN NAND3X2 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 1.300000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.602000 0.300000 0.698000 0.490000 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.782000 0.433000 0.907000 0.588000 ;
        RECT 0.782000 0.493000 0.923000 0.588000 ;
        RECT 0.377000 0.514000 0.473000 0.604000 ;
        RECT 0.782000 0.433000 0.868000 0.604000 ;
        RECT 0.377000 0.549000 0.868000 0.604000 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.087000 0.460000 0.183000 0.573000 ;
        RECT 1.016000 0.573000 1.111000 0.706000 ;
        RECT 0.087000 0.439000 0.167000 0.573000 ;
        RECT 1.031000 0.573000 1.096000 0.881000 ;
        RECT 0.118000 0.460000 0.183000 0.881000 ;
        RECT 0.118000 0.826000 1.096000 0.881000 ;
        RECT 0.060000 0.439000 0.167000 0.494000 ;
        RECT 0.118000 0.439000 0.167000 0.881000 ;
        END
    END C
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 1.300000 1.280000 ;
        RECT 0.499000 0.952000 0.595000 1.280000 ;
        RECT 0.108000 0.952000 0.204000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 1.300000 0.080000 ;
        RECT 1.137000 -0.080000 1.232000 0.122000 ;
        RECT 0.068000 -0.080000 0.163000 0.122000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.691000 0.689000 0.786000 0.770000 ;
        RECT 0.602000 0.164000 0.698000 0.245000 ;
        RECT 0.300000 0.689000 0.432000 0.770000 ;
        RECT 0.682000 0.689000 0.786000 0.761000 ;
        RECT 0.248000 0.689000 0.432000 0.761000 ;
        RECT 0.300000 0.700000 0.518000 0.770000 ;
        RECT 0.248000 0.190000 0.312000 0.761000 ;
        RECT 0.248000 0.700000 0.518000 0.761000 ;
        RECT 0.248000 0.706000 0.786000 0.761000 ;
        RECT 0.248000 0.190000 0.698000 0.245000 ;
        RECT 0.300000 0.190000 0.312000 0.770000 ;
        END
    END Y
END NAND3X2

MACRO NAND2BX4
    CLASS CORE ;
    FOREIGN NAND2BX4 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 1.400000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN AN
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.045000 0.481000 0.135000 0.633000 ;
        END
    END AN
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.818000 0.568000 0.985000 0.662000 ;
        RECT 0.334000 0.568000 0.424000 0.662000 ;
        RECT 0.334000 0.573000 0.480000 0.662000 ;
        RECT 0.334000 0.607000 0.985000 0.662000 ;
        END
    END B
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 1.400000 1.280000 ;
        RECT 0.905000 0.871000 0.996000 1.280000 ;
        RECT 1.246000 0.871000 1.336000 1.280000 ;
        RECT 0.566000 0.871000 0.656000 1.280000 ;
        RECT 0.227000 0.883000 0.317000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 1.400000 0.080000 ;
        RECT 0.923000 -0.080000 1.013000 0.254000 ;
        RECT 0.249000 -0.080000 0.339000 0.122000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.262000 0.245000 1.363000 0.633000 ;
        RECT 1.267000 0.245000 1.358000 0.798000 ;
        RECT 0.583000 0.283000 0.673000 0.399000 ;
        RECT 0.396000 0.717000 1.358000 0.798000 ;
        RECT 0.583000 0.327000 1.363000 0.399000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 0.581000 0.457000 0.671000 0.552000 ;
        RECT 0.048000 0.717000 0.138000 0.798000 ;
        RECT 0.048000 0.279000 0.138000 0.360000 ;
        RECT 1.140000 0.457000 1.201000 0.649000 ;
        RECT 0.199000 0.305000 0.260000 0.771000 ;
        RECT 0.581000 0.457000 1.201000 0.512000 ;
        RECT 0.260000 0.457000 0.581000 0.512000 ;
        RECT 0.048000 0.305000 0.260000 0.360000 ;
        RECT 0.048000 0.717000 0.260000 0.771000 ;
    END
END NAND2BX4

MACRO NAND2BX2
    CLASS CORE ;
    FOREIGN NAND2BX2 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 1.100000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN AN
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.047000 0.452000 0.142000 0.627000 ;
        END
    END AN
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.853000 0.549000 0.939000 0.636000 ;
        RECT 0.372000 0.560000 0.467000 0.640000 ;
        RECT 0.372000 0.573000 0.939000 0.627000 ;
        END
    END B
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.353000 1.078000 1.050000 1.280000 ;
        RECT 0.000000 1.120000 1.100000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 1.100000 0.080000 ;
        RECT 0.233000 -0.080000 0.328000 0.122000 ;
        RECT 0.956000 -0.080000 1.050000 0.278000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.800000 0.690000 0.894000 0.771000 ;
        RECT 0.600000 0.290000 0.694000 0.371000 ;
        RECT 0.444000 0.702000 0.539000 0.783000 ;
        RECT 0.772000 0.700000 1.067000 0.770000 ;
        RECT 0.444000 0.702000 0.610000 0.770000 ;
        RECT 0.812000 0.361000 0.878000 0.457000 ;
        RECT 1.003000 0.402000 1.067000 0.770000 ;
        RECT 0.812000 0.317000 0.876000 0.457000 ;
        RECT 0.812000 0.402000 1.067000 0.457000 ;
        RECT 0.444000 0.715000 1.067000 0.770000 ;
        RECT 0.600000 0.317000 0.876000 0.371000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 0.050000 0.279000 0.144000 0.368000 ;
        RECT 0.639000 0.433000 0.733000 0.514000 ;
        RECT 0.050000 0.702000 0.144000 0.783000 ;
        RECT 0.049000 0.292000 0.144000 0.368000 ;
        RECT 0.208000 0.311000 0.272000 0.757000 ;
        RECT 0.049000 0.311000 0.272000 0.368000 ;
        RECT 0.272000 0.446000 0.639000 0.501000 ;
        RECT 0.050000 0.702000 0.272000 0.757000 ;
    END
END NAND2BX2

MACRO NAND2X4
    CLASS CORE ;
    FOREIGN NAND2X4 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 1.300000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.968000 0.467000 1.089000 0.573000 ;
        RECT 0.605000 0.439000 0.695000 0.521000 ;
        RECT 0.431000 0.471000 0.526000 0.552000 ;
        RECT 0.446000 0.467000 0.526000 0.552000 ;
        RECT 1.024000 0.467000 1.089000 0.652000 ;
        RECT 0.446000 0.467000 1.089000 0.521000 ;
        RECT 0.431000 0.471000 1.089000 0.521000 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.184000 0.573000 0.311000 0.662000 ;
        RECT 0.764000 0.576000 0.860000 0.657000 ;
        RECT 0.169000 0.573000 0.311000 0.654000 ;
        RECT 0.764000 0.576000 0.844000 0.662000 ;
        RECT 0.184000 0.607000 0.844000 0.662000 ;
        RECT 0.184000 0.607000 0.860000 0.657000 ;
        END
    END B
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 1.300000 1.280000 ;
        RECT 1.131000 0.871000 1.227000 1.280000 ;
        RECT 0.771000 0.871000 0.867000 1.280000 ;
        RECT 0.411000 0.871000 0.506000 1.280000 ;
        RECT 0.051000 0.871000 0.146000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 1.300000 0.080000 ;
        RECT 0.794000 -0.080000 0.889000 0.237000 ;
        RECT 0.079000 -0.080000 0.174000 0.122000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.154000 0.245000 1.261000 0.633000 ;
        RECT 0.433000 0.283000 0.529000 0.379000 ;
        RECT 1.154000 0.245000 1.249000 0.798000 ;
        RECT 0.231000 0.717000 1.249000 0.798000 ;
        RECT 0.433000 0.307000 1.261000 0.379000 ;
        END
    END Y
END NAND2X4

MACRO NAND2X2
    CLASS CORE ;
    FOREIGN NAND2X2 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 0.900000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.398000 0.400000 0.551000 0.520000 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.668000 0.558000 0.731000 0.645000 ;
        RECT 0.200000 0.573000 0.301000 0.632000 ;
        RECT 0.200000 0.577000 0.731000 0.632000 ;
        RECT 0.185000 0.573000 0.301000 0.627000 ;
        RECT 0.185000 0.577000 0.731000 0.627000 ;
        END
    END B
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.210000 1.078000 0.851000 1.280000 ;
        RECT 0.000000 1.120000 0.900000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 0.900000 0.080000 ;
        RECT 0.758000 -0.080000 0.851000 0.289000 ;
        RECT 0.049000 -0.080000 0.142000 0.122000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.409000 0.223000 0.502000 0.304000 ;
        RECT 0.779000 0.704000 0.858000 0.770000 ;
        RECT 0.795000 0.402000 0.858000 0.770000 ;
        RECT 0.618000 0.249000 0.680000 0.457000 ;
        RECT 0.599000 0.249000 0.680000 0.306000 ;
        RECT 0.618000 0.402000 0.858000 0.457000 ;
        RECT 0.409000 0.249000 0.680000 0.304000 ;
        RECT 0.251000 0.704000 0.858000 0.758000 ;
        END
    END Y
END NAND2X2

MACRO MXI4X2
    CLASS CORE ;
    FOREIGN MXI4X2 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 4.200000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.037000 0.526000 0.209000 0.633000 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.862000 0.450000 0.969000 0.527000 ;
        RECT 0.908000 0.306000 0.969000 0.527000 ;
        RECT 0.908000 0.306000 0.993000 0.361000 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 2.205000 0.474000 2.292000 0.561000 ;
        RECT 2.233000 0.300000 2.413000 0.367000 ;
        RECT 2.231000 0.306000 2.413000 0.367000 ;
        RECT 2.231000 0.306000 2.292000 0.561000 ;
        RECT 2.233000 0.300000 2.292000 0.561000 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.437000 0.302000 1.548000 0.533000 ;
        END
    END D
    PIN S0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.053000 0.433000 1.188000 0.567000 ;
        END
    END S0
    PIN S1
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 3.187000 0.433000 3.371000 0.524000 ;
        END
    END S1
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 4.200000 1.280000 ;
        RECT 3.810000 1.078000 3.900000 1.280000 ;
        RECT 3.344000 1.078000 3.434000 1.280000 ;
        RECT 2.270000 1.078000 2.360000 1.280000 ;
        RECT 1.379000 0.954000 1.469000 1.280000 ;
        RECT 0.952000 0.954000 1.042000 1.280000 ;
        RECT 0.061000 0.745000 0.151000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 4.200000 0.080000 ;
        RECT 3.834000 -0.080000 3.924000 0.122000 ;
        RECT 3.378000 -0.080000 3.468000 0.122000 ;
        RECT 2.270000 -0.080000 2.360000 0.217000 ;
        RECT 1.432000 -0.080000 1.522000 0.217000 ;
        RECT 0.952000 -0.080000 1.042000 0.220000 ;
        RECT 0.061000 -0.080000 0.151000 0.329000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 3.887000 0.665000 4.148000 0.767000 ;
        RECT 4.049000 0.665000 4.148000 1.007000 ;
        RECT 4.052000 0.183000 4.148000 0.376000 ;
        RECT 4.082000 0.627000 4.148000 1.007000 ;
        RECT 4.087000 0.183000 4.148000 1.007000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 3.177000 0.637000 3.273000 0.735000 ;
        RECT 3.011000 0.445000 3.106000 0.545000 ;
        RECT 3.448000 0.761000 3.639000 0.854000 ;
        RECT 2.873000 0.767000 2.986000 0.854000 ;
        RECT 2.873000 0.287000 2.955000 0.374000 ;
        RECT 3.914000 0.496000 4.004000 0.577000 ;
        RECT 3.590000 0.514000 3.680000 0.595000 ;
        RECT 2.693000 0.796000 2.780000 0.877000 ;
        RECT 2.678000 0.262000 2.768000 0.343000 ;
        RECT 1.851000 0.252000 1.990000 0.333000 ;
        RECT 1.649000 0.252000 1.739000 0.333000 ;
        RECT 0.420000 0.237000 0.570000 0.318000 ;
        RECT 0.711000 0.260000 0.801000 0.340000 ;
        RECT 3.605000 0.514000 3.680000 0.596000 ;
        RECT 3.914000 0.198000 3.975000 0.577000 ;
        RECT 3.716000 0.542000 3.777000 1.008000 ;
        RECT 3.448000 0.313000 3.509000 0.854000 ;
        RECT 3.249000 0.163000 3.310000 0.252000 ;
        RECT 3.045000 0.313000 3.106000 0.692000 ;
        RECT 2.873000 0.287000 2.934000 0.854000 ;
        RECT 2.707000 0.163000 2.768000 0.343000 ;
        RECT 2.693000 0.262000 2.754000 0.877000 ;
        RECT 2.528000 0.177000 2.589000 0.877000 ;
        RECT 2.401000 0.495000 2.462000 0.898000 ;
        RECT 2.067000 0.252000 2.128000 0.776000 ;
        RECT 1.929000 0.252000 1.990000 0.898000 ;
        RECT 1.791000 0.436000 1.852000 0.774000 ;
        RECT 1.678000 0.252000 1.739000 0.490000 ;
        RECT 1.653000 0.546000 1.714000 0.664000 ;
        RECT 1.584000 0.830000 1.645000 1.008000 ;
        RECT 1.269000 0.287000 1.330000 0.744000 ;
        RECT 0.866000 0.595000 0.927000 0.744000 ;
        RECT 0.711000 0.260000 0.772000 0.439000 ;
        RECT 0.696000 0.510000 0.757000 0.650000 ;
        RECT 0.558000 0.385000 0.619000 0.760000 ;
        RECT 0.420000 0.237000 0.481000 0.885000 ;
        RECT 0.282000 0.263000 0.343000 0.817000 ;
        RECT 3.448000 0.313000 3.717000 0.368000 ;
        RECT 3.045000 0.637000 3.273000 0.692000 ;
        RECT 3.045000 0.313000 3.166000 0.368000 ;
        RECT 2.873000 0.799000 3.639000 0.854000 ;
        RECT 2.707000 0.163000 3.310000 0.218000 ;
        RECT 2.477000 0.177000 2.589000 0.232000 ;
        RECT 1.787000 0.843000 2.462000 0.898000 ;
        RECT 1.586000 0.719000 1.852000 0.774000 ;
        RECT 1.169000 0.287000 1.330000 0.342000 ;
        RECT 0.866000 0.689000 1.330000 0.744000 ;
        RECT 0.696000 0.595000 0.927000 0.650000 ;
        RECT 0.558000 0.705000 0.782000 0.760000 ;
        RECT 0.420000 0.830000 1.645000 0.885000 ;
        RECT 3.605000 0.542000 3.777000 0.596000 ;
        RECT 3.249000 0.198000 3.975000 0.252000 ;
        RECT 1.678000 0.436000 1.852000 0.490000 ;
        RECT 1.584000 0.954000 3.777000 1.008000 ;
        RECT 1.269000 0.610000 1.714000 0.664000 ;
        RECT 0.558000 0.385000 0.772000 0.439000 ;
        RECT 3.590000 0.542000 3.777000 0.595000 ;
        RECT 2.707000 0.163000 2.754000 0.877000 ;
    END
END MXI4X2

MACRO MXI2X4
    CLASS CORE ;
    FOREIGN MXI2X4 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 2.500000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.152000 0.526000 0.406000 0.607000 ;
        RECT 0.237000 0.526000 0.299000 0.627000 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 2.002000 0.514000 2.189000 0.633000 ;
        END
    END B
    PIN S0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.602000 0.954000 1.694000 1.035000 ;
        RECT 1.466000 0.967000 1.694000 1.035000 ;
        RECT 0.564000 0.943000 0.626000 1.035000 ;
        RECT 0.564000 0.980000 1.694000 1.035000 ;
        END
    END S0
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 2.500000 1.280000 ;
        RECT 2.359000 0.979000 2.451000 1.280000 ;
        RECT 1.979000 0.896000 2.071000 1.280000 ;
        RECT 0.054000 0.982000 0.146000 1.280000 ;
        RECT 0.421000 0.979000 0.483000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 2.500000 0.080000 ;
        RECT 2.359000 -0.080000 2.451000 0.235000 ;
        RECT 1.986000 -0.080000 2.078000 0.122000 ;
        RECT 0.407000 -0.080000 0.499000 0.235000 ;
        RECT 0.054000 -0.080000 0.146000 0.240000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.109000 0.167000 1.212000 0.500000 ;
        RECT 1.518000 0.171000 1.604000 0.262000 ;
        RECT 1.109000 0.171000 1.215000 0.255000 ;
        RECT 0.736000 0.171000 0.828000 0.252000 ;
        RECT 1.013000 0.833000 1.155000 0.908000 ;
        RECT 1.093000 0.439000 1.155000 0.908000 ;
        RECT 1.093000 0.439000 1.212000 0.500000 ;
        RECT 0.736000 0.171000 1.604000 0.226000 ;
        RECT 0.694000 0.854000 1.527000 0.908000 ;
        RECT 1.109000 0.167000 1.155000 0.908000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 1.792000 0.662000 1.893000 0.764000 ;
        RECT 2.179000 0.705000 2.271000 0.865000 ;
        RECT 0.874000 0.657000 0.966000 0.751000 ;
        RECT 0.233000 0.336000 0.325000 0.449000 ;
        RECT 0.233000 0.699000 0.325000 0.786000 ;
        RECT 2.181000 0.336000 2.273000 0.417000 ;
        RECT 1.243000 0.679000 1.335000 0.760000 ;
        RECT 0.908000 0.336000 1.000000 0.417000 ;
        RECT 1.602000 0.710000 1.694000 0.790000 ;
        RECT 2.196000 0.336000 2.273000 0.418000 ;
        RECT 0.248000 0.696000 0.325000 0.786000 ;
        RECT 2.179000 0.336000 2.273000 0.404000 ;
        RECT 2.344000 0.363000 2.407000 0.760000 ;
        RECT 2.179000 0.221000 2.242000 0.404000 ;
        RECT 1.792000 0.336000 1.855000 0.764000 ;
        RECT 1.339000 0.349000 1.402000 0.733000 ;
        RECT 1.668000 0.221000 1.730000 0.404000 ;
        RECT 0.813000 0.362000 0.875000 0.449000 ;
        RECT 0.499000 0.394000 0.561000 0.754000 ;
        RECT 2.181000 0.221000 2.242000 0.417000 ;
        RECT 0.248000 0.696000 0.561000 0.754000 ;
        RECT 2.196000 0.363000 2.407000 0.418000 ;
        RECT 2.179000 0.705000 2.407000 0.760000 ;
        RECT 1.668000 0.221000 2.242000 0.276000 ;
        RECT 1.339000 0.349000 1.730000 0.404000 ;
        RECT 0.813000 0.362000 1.000000 0.417000 ;
        RECT 0.248000 0.696000 0.966000 0.751000 ;
        RECT 0.233000 0.699000 0.561000 0.754000 ;
        RECT 0.233000 0.394000 0.875000 0.449000 ;
        RECT 2.181000 0.363000 2.407000 0.417000 ;
        RECT 1.602000 0.710000 1.893000 0.764000 ;
        RECT 1.243000 0.679000 1.402000 0.733000 ;
        RECT 0.233000 0.699000 0.966000 0.751000 ;
        RECT 2.196000 0.221000 2.242000 0.418000 ;
    END
END MXI2X4

MACRO MXI2X2
    CLASS CORE ;
    FOREIGN MXI2X2 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 1.400000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.252000 0.433000 1.363000 0.576000 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.387000 0.506000 0.493000 0.633000 ;
        END
    END B
    PIN S0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.179000 0.656000 0.313000 0.767000 ;
        END
    END S0
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 1.400000 1.280000 ;
        RECT 0.286000 0.853000 0.377000 1.280000 ;
        RECT 1.262000 0.757000 1.352000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 1.400000 0.080000 ;
        RECT 1.262000 -0.080000 1.352000 0.122000 ;
        RECT 0.369000 -0.080000 0.459000 0.261000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.716000 0.833000 0.838000 1.005000 ;
        RECT 0.883000 0.293000 0.944000 0.888000 ;
        RECT 0.716000 0.833000 0.944000 0.888000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 1.025000 0.736000 1.115000 0.960000 ;
        RECT 0.554000 0.517000 0.696000 0.607000 ;
        RECT 0.493000 0.708000 0.583000 1.013000 ;
        RECT 0.167000 0.257000 0.257000 0.348000 ;
        RECT 0.677000 0.326000 0.822000 0.407000 ;
        RECT 0.048000 0.836000 0.138000 0.917000 ;
        RECT 1.128000 0.336000 1.189000 0.790000 ;
        RECT 1.005000 0.163000 1.066000 0.571000 ;
        RECT 0.761000 0.326000 0.822000 0.763000 ;
        RECT 0.554000 0.163000 0.615000 0.607000 ;
        RECT 0.196000 0.257000 0.257000 0.442000 ;
        RECT 0.048000 0.293000 0.109000 0.917000 ;
        RECT 0.554000 0.163000 1.066000 0.218000 ;
        RECT 0.493000 0.708000 0.822000 0.763000 ;
        RECT 0.196000 0.387000 0.615000 0.442000 ;
        RECT 0.048000 0.293000 0.257000 0.348000 ;
        RECT 1.025000 0.736000 1.189000 0.790000 ;
    END
END MXI2X2

MACRO MX2X4
    CLASS CORE ;
    FOREIGN MX2X4 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 1.800000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.118000 0.433000 1.261000 0.533000 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.235000 0.421000 0.413000 0.512000 ;
        RECT 0.218000 0.433000 0.413000 0.512000 ;
        END
    END B
    PIN S0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.170000 0.677000 0.266000 0.767000 ;
        RECT 0.170000 0.700000 0.502000 0.767000 ;
        END
    END S0
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 1.800000 1.280000 ;
        RECT 1.227000 0.986000 1.320000 1.280000 ;
        RECT 0.262000 0.855000 0.355000 1.280000 ;
        RECT 1.653000 1.078000 1.745000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 1.800000 0.080000 ;
        RECT 1.655000 -0.080000 1.748000 0.211000 ;
        RECT 1.279000 -0.080000 1.372000 0.211000 ;
        RECT 0.305000 -0.080000 0.398000 0.352000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.478000 0.167000 1.582000 0.798000 ;
        RECT 1.424000 0.707000 1.582000 0.798000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 0.494000 0.475000 0.642000 0.557000 ;
        RECT 1.651000 0.495000 1.744000 0.576000 ;
        RECT 1.001000 0.707000 1.094000 0.788000 ;
        RECT 0.712000 0.833000 0.919000 0.914000 ;
        RECT 0.620000 0.290000 0.772000 0.371000 ;
        RECT 0.475000 0.837000 0.567000 0.918000 ;
        RECT 0.045000 0.840000 0.147000 0.921000 ;
        RECT 0.045000 0.293000 0.147000 0.374000 ;
        RECT 1.666000 0.495000 1.729000 0.914000 ;
        RECT 1.324000 0.313000 1.387000 0.651000 ;
        RECT 1.031000 0.596000 1.094000 0.788000 ;
        RECT 0.982000 0.161000 1.045000 0.507000 ;
        RECT 0.856000 0.290000 0.919000 0.914000 ;
        RECT 0.709000 0.290000 0.772000 0.758000 ;
        RECT 0.585000 0.704000 0.648000 0.892000 ;
        RECT 0.045000 0.293000 0.108000 0.921000 ;
        RECT 0.494000 0.161000 0.556000 0.621000 ;
        RECT 1.107000 0.313000 1.387000 0.368000 ;
        RECT 1.031000 0.596000 1.387000 0.651000 ;
        RECT 0.475000 0.837000 0.648000 0.892000 ;
        RECT 0.712000 0.860000 1.729000 0.914000 ;
        RECT 0.585000 0.704000 0.772000 0.758000 ;
        RECT 0.494000 0.161000 1.045000 0.215000 ;
        RECT 0.045000 0.567000 0.556000 0.621000 ;
    END
END MX2X4

MACRO MX2X2
    CLASS CORE ;
    FOREIGN MX2X2 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 1.600000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.160000 0.306000 1.222000 0.575000 ;
        RECT 1.160000 0.306000 1.285000 0.367000 ;
        RECT 1.160000 0.306000 1.364000 0.361000 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.215000 0.526000 0.387000 0.633000 ;
        END
    END B
    PIN S0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.210000 0.714000 0.302000 0.795000 ;
        RECT 0.225000 0.706000 0.302000 0.795000 ;
        RECT 0.225000 0.706000 0.475000 0.761000 ;
        END
    END S0
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 1.600000 1.280000 ;
        RECT 1.231000 1.078000 1.323000 1.280000 ;
        RECT 0.315000 0.890000 0.407000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 1.600000 0.080000 ;
        RECT 1.244000 -0.080000 1.336000 0.223000 ;
        RECT 0.315000 -0.080000 0.407000 0.296000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.446000 0.700000 1.556000 0.977000 ;
        RECT 1.461000 0.194000 1.556000 0.395000 ;
        RECT 1.480000 0.194000 1.556000 0.439000 ;
        RECT 1.494000 0.194000 1.556000 0.977000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 1.323000 0.485000 1.415000 0.595000 ;
        RECT 0.770000 0.836000 0.941000 0.917000 ;
        RECT 0.752000 0.240000 0.843000 0.321000 ;
        RECT 0.054000 0.858000 0.145000 0.939000 ;
        RECT 0.048000 0.348000 0.140000 0.429000 ;
        RECT 1.323000 0.485000 1.385000 0.994000 ;
        RECT 0.879000 0.267000 0.941000 0.994000 ;
        RECT 0.739000 0.396000 0.801000 0.761000 ;
        RECT 0.605000 0.190000 0.667000 0.451000 ;
        RECT 0.599000 0.520000 0.661000 0.606000 ;
        RECT 0.580000 0.706000 0.642000 0.915000 ;
        RECT 0.465000 0.370000 0.527000 0.575000 ;
        RECT 0.063000 0.348000 0.125000 0.939000 ;
        RECT 1.020000 0.279000 1.081000 0.858000 ;
        RECT 0.879000 0.939000 1.385000 0.994000 ;
        RECT 0.605000 0.396000 0.801000 0.451000 ;
        RECT 0.580000 0.706000 0.801000 0.761000 ;
        RECT 0.547000 0.190000 0.667000 0.245000 ;
        RECT 0.465000 0.520000 0.661000 0.575000 ;
        RECT 0.145000 0.370000 0.527000 0.425000 ;
        RECT 0.140000 0.370000 0.465000 0.425000 ;
        RECT 0.048000 0.370000 0.145000 0.425000 ;
        RECT 0.752000 0.267000 0.941000 0.321000 ;
    END
END MX2X2

MACRO INVX8
    CLASS CORE ;
    FOREIGN INVX8 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 1.100000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.150000 0.487000 0.376000 0.633000 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.828000 1.078000 1.050000 1.280000 ;
        RECT 0.000000 1.120000 1.100000 1.280000 ;
        RECT 0.828000 0.917000 0.922000 1.280000 ;
        RECT 0.438000 0.917000 0.532000 1.280000 ;
        RECT 0.050000 0.917000 0.144000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.818000 -0.080000 1.043000 0.122000 ;
        RECT 0.000000 -0.080000 1.100000 0.080000 ;
        RECT 0.061000 -0.080000 0.156000 0.122000 ;
        RECT 0.439000 -0.080000 0.533000 0.214000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.610000 0.419000 1.040000 0.767000 ;
        RECT 0.610000 0.361000 0.878000 0.767000 ;
        RECT 0.610000 0.361000 0.857000 0.780000 ;
        RECT 0.610000 0.307000 0.811000 0.812000 ;
        RECT 0.589000 0.307000 0.811000 0.433000 ;
        RECT 0.217000 0.698000 0.811000 0.812000 ;
        RECT 0.217000 0.307000 0.811000 0.421000 ;
        RECT 0.217000 0.698000 0.857000 0.780000 ;
        RECT 0.589000 0.361000 0.878000 0.433000 ;
        RECT 0.217000 0.698000 1.040000 0.767000 ;
        RECT 0.217000 0.361000 0.878000 0.421000 ;
        END
    END Y
END INVX8

MACRO INVX4
    CLASS CORE ;
    FOREIGN INVX4 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 0.700000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.037000 0.446000 0.138000 0.633000 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 0.700000 1.280000 ;
        RECT 0.452000 0.720000 0.542000 1.280000 ;
        RECT 0.048000 0.720000 0.138000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 0.700000 0.080000 ;
        RECT 0.452000 -0.080000 0.542000 0.372000 ;
        RECT 0.048000 -0.080000 0.138000 0.372000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.212000 0.433000 0.341000 0.767000 ;
        RECT 0.251000 0.194000 0.341000 1.010000 ;
        END
    END Y
END INVX4

MACRO INVX3
    CLASS CORE ;
    FOREIGN INVX3 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 0.700000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.037000 0.493000 0.266000 0.633000 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 0.700000 1.280000 ;
        RECT 0.251000 1.078000 0.341000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 0.700000 0.080000 ;
        RECT 0.251000 -0.080000 0.341000 0.122000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.387000 0.700000 0.489000 0.900000 ;
        RECT 0.399000 0.295000 0.489000 0.913000 ;
        RECT 0.049000 0.720000 0.139000 0.913000 ;
        RECT 0.049000 0.215000 0.139000 0.408000 ;
        RECT 0.049000 0.773000 0.489000 0.854000 ;
        RECT 0.049000 0.295000 0.489000 0.376000 ;
        END
    END Y
END INVX3

MACRO INVX2
    CLASS CORE ;
    FOREIGN INVX2 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 0.600000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.150000 0.433000 0.395000 0.574000 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 0.600000 1.280000 ;
        RECT 0.394000 1.078000 0.497000 1.280000 ;
        RECT 0.395000 1.064000 0.495000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 0.600000 0.080000 ;
        RECT 0.164000 -0.080000 0.267000 0.361000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.442000 0.183000 0.558000 0.376000 ;
        RECT 0.224000 0.661000 0.327000 0.854000 ;
        RECT 0.465000 0.627000 0.558000 0.715000 ;
        RECT 0.488000 0.183000 0.558000 0.715000 ;
        RECT 0.224000 0.661000 0.558000 0.715000 ;
        END
    END Y
END INVX2

MACRO DFFX2
    CLASS CORE ;
    FOREIGN DFFX2 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 3.700000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER Metal1 ;
        RECT 0.214000 0.505000 0.315000 0.633000 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.390000 0.335000 0.487000 0.494000 ;
        RECT 0.354000 0.335000 0.487000 0.415000 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 2.995000 0.167000 3.086000 0.248000 ;
        RECT 2.888000 0.683000 2.979000 0.764000 ;
        RECT 2.995000 0.167000 3.071000 0.257000 ;
        RECT 2.888000 0.567000 2.958000 0.764000 ;
        RECT 2.856000 0.567000 2.958000 0.633000 ;
        RECT 2.839000 0.202000 2.900000 0.621000 ;
        RECT 2.839000 0.202000 3.071000 0.257000 ;
        RECT 2.839000 0.567000 2.958000 0.621000 ;
        RECT 2.856000 0.202000 2.888000 0.633000 ;
        RECT 2.888000 0.202000 2.900000 0.764000 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 3.385000 0.323000 3.466000 0.439000 ;
        RECT 3.358000 0.323000 3.466000 0.404000 ;
        RECT 3.300000 0.738000 3.390000 0.819000 ;
        RECT 3.405000 0.323000 3.466000 0.793000 ;
        RECT 3.300000 0.738000 3.466000 0.793000 ;
        END
    END QN
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 2.186000 1.078000 2.654000 1.280000 ;
        RECT 0.000000 1.120000 3.700000 1.280000 ;
        RECT 3.449000 1.078000 3.540000 1.280000 ;
        RECT 3.091000 1.078000 3.182000 1.280000 ;
        RECT 0.296000 1.065000 0.387000 1.280000 ;
        RECT 1.482000 1.078000 1.572000 1.280000 ;
        RECT 1.119000 1.078000 1.209000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 3.700000 0.080000 ;
        RECT 3.508000 -0.080000 3.599000 0.122000 ;
        RECT 3.209000 -0.080000 3.300000 0.122000 ;
        RECT 2.258000 -0.080000 2.349000 0.287000 ;
        RECT 1.560000 -0.080000 1.651000 0.329000 ;
        RECT 0.982000 -0.080000 1.073000 0.287000 ;
        RECT 0.203000 -0.080000 0.294000 0.122000 ;
        RECT 2.782000 -0.080000 2.872000 0.122000 ;
        END
    END VSS
    OBS
        LAYER Metal1 ;
        RECT 0.243000 0.719000 0.350000 0.913000 ;
        RECT 2.472000 0.275000 2.563000 0.427000 ;
        RECT 2.888000 0.951000 2.979000 1.040000 ;
        RECT 3.244000 0.957000 3.334000 1.038000 ;
        RECT 2.320000 0.800000 2.411000 0.881000 ;
        RECT 1.917000 0.250000 2.008000 0.331000 ;
        RECT 1.858000 0.671000 1.949000 0.752000 ;
        RECT 1.352000 0.263000 1.454000 0.344000 ;
        RECT 1.332000 0.625000 1.423000 0.706000 ;
        RECT 0.957000 0.517000 1.251000 0.598000 ;
        RECT 0.619000 0.193000 0.710000 0.274000 ;
        RECT 0.558000 0.329000 0.649000 0.410000 ;
        RECT 0.048000 0.319000 0.152000 0.400000 ;
        RECT 2.432000 0.560000 2.523000 0.640000 ;
        RECT 3.244000 0.951000 3.320000 1.038000 ;
        RECT 0.884000 0.926000 0.960000 1.006000 ;
        RECT 2.320000 0.800000 2.663000 0.874000 ;
        RECT 3.175000 0.368000 3.237000 1.006000 ;
        RECT 2.888000 0.929000 2.950000 1.040000 ;
        RECT 2.601000 0.423000 2.663000 0.874000 ;
        RECT 2.501000 0.275000 2.563000 0.477000 ;
        RECT 2.126000 0.573000 2.188000 0.752000 ;
        RECT 1.863000 0.425000 1.925000 0.752000 ;
        RECT 1.628000 0.698000 1.690000 1.008000 ;
        RECT 1.352000 0.150000 1.414000 0.706000 ;
        RECT 1.189000 0.226000 1.251000 0.598000 ;
        RECT 0.898000 0.926000 0.960000 1.008000 ;
        RECT 0.881000 0.926000 0.960000 0.988000 ;
        RECT 0.834000 0.368000 0.896000 0.857000 ;
        RECT 0.731000 0.219000 0.793000 0.425000 ;
        RECT 0.711000 0.671000 0.773000 0.981000 ;
        RECT 0.467000 0.858000 0.529000 0.981000 ;
        RECT 3.053000 0.544000 3.114000 0.874000 ;
        RECT 2.320000 0.800000 2.381000 0.943000 ;
        RECT 2.109000 0.276000 2.170000 0.427000 ;
        RECT 1.849000 0.819000 1.910000 1.018000 ;
        RECT 1.503000 0.535000 1.564000 0.899000 ;
        RECT 1.192000 0.540000 1.253000 0.899000 ;
        RECT 0.573000 0.329000 0.634000 0.726000 ;
        RECT 0.091000 0.319000 0.152000 0.788000 ;
        RECT 1.192000 0.226000 1.251000 0.899000 ;
        RECT 0.957000 0.540000 1.253000 0.598000 ;
        RECT 0.731000 0.368000 0.896000 0.425000 ;
        RECT 2.995000 0.368000 3.237000 0.423000 ;
        RECT 2.979000 0.951000 3.320000 1.006000 ;
        RECT 2.888000 0.951000 3.237000 1.006000 ;
        RECT 2.320000 0.819000 3.114000 0.874000 ;
        RECT 1.917000 0.276000 2.170000 0.331000 ;
        RECT 1.849000 0.888000 2.381000 0.943000 ;
        RECT 1.476000 0.425000 1.925000 0.480000 ;
        RECT 1.317000 0.150000 1.414000 0.205000 ;
        RECT 1.192000 0.844000 1.564000 0.899000 ;
        RECT 0.731000 0.370000 1.116000 0.425000 ;
        RECT 0.619000 0.219000 0.793000 0.274000 ;
        RECT 0.573000 0.671000 0.773000 0.726000 ;
        RECT 0.467000 0.926000 0.960000 0.981000 ;
        RECT 0.243000 0.858000 0.529000 0.913000 ;
        RECT 0.091000 0.733000 0.350000 0.788000 ;
        RECT 2.573000 0.929000 2.950000 0.983000 ;
        RECT 2.501000 0.423000 2.663000 0.477000 ;
        RECT 2.126000 0.573000 2.523000 0.627000 ;
        RECT 2.109000 0.373000 2.563000 0.427000 ;
        RECT 1.628000 0.698000 2.188000 0.752000 ;
        RECT 1.503000 0.535000 1.765000 0.589000 ;
        RECT 0.898000 0.954000 1.690000 1.008000 ;
        RECT 0.884000 0.954000 1.690000 1.006000 ;
    END
END DFFX2

MACRO BUFX8
    CLASS CORE ;
    FOREIGN BUFX8 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 1.600000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.154000 0.474000 0.372000 0.555000 ;
        RECT 0.236000 0.439000 0.298000 0.555000 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 1.600000 1.280000 ;
        RECT 1.104000 0.877000 1.196000 1.280000 ;
        RECT 0.070000 0.897000 0.162000 1.280000 ;
        RECT 0.760000 0.877000 0.851000 1.280000 ;
        RECT 0.415000 0.897000 0.506000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 1.600000 0.080000 ;
        RECT 1.126000 -0.080000 1.218000 0.211000 ;
        RECT 0.781000 -0.080000 0.873000 0.211000 ;
        RECT 0.436000 -0.080000 0.528000 0.198000 ;
        RECT 0.048000 -0.080000 0.140000 0.211000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.947000 0.433000 1.364000 0.767000 ;
        RECT 0.947000 0.433000 1.220000 0.774000 ;
        RECT 0.947000 0.307000 1.131000 0.774000 ;
        RECT 0.927000 0.626000 1.220000 0.774000 ;
        RECT 0.927000 0.626000 1.364000 0.767000 ;
        RECT 0.927000 0.307000 1.131000 0.440000 ;
        RECT 0.609000 0.307000 1.131000 0.421000 ;
        RECT 0.587000 0.660000 1.220000 0.774000 ;
        RECT 0.587000 0.660000 1.364000 0.767000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 0.434000 0.274000 0.525000 0.738000 ;
        RECT 0.434000 0.519000 0.865000 0.600000 ;
        RECT 0.242000 0.657000 0.525000 0.738000 ;
        RECT 0.242000 0.274000 0.525000 0.355000 ;
    END
END BUFX8

MACRO BUFX4
    CLASS CORE ;
    FOREIGN BUFX4 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 0.900000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.038000 0.433000 0.218000 0.570000 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 0.900000 1.280000 ;
        RECT 0.671000 0.953000 0.764000 1.280000 ;
        RECT 0.256000 0.953000 0.349000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 0.900000 0.080000 ;
        RECT 0.671000 -0.080000 0.764000 0.122000 ;
        RECT 0.256000 -0.080000 0.349000 0.122000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.464000 0.652000 0.600000 0.767000 ;
        RECT 0.464000 0.300000 0.682000 0.412000 ;
        RECT 0.578000 0.300000 0.682000 0.733000 ;
        RECT 0.464000 0.652000 0.556000 0.957000 ;
        RECT 0.464000 0.219000 0.556000 0.412000 ;
        RECT 0.464000 0.652000 0.682000 0.733000 ;
        RECT 0.578000 0.300000 0.600000 0.767000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 0.284000 0.477000 0.515000 0.585000 ;
        RECT 0.049000 0.652000 0.142000 0.957000 ;
        RECT 0.049000 0.186000 0.142000 0.379000 ;
        RECT 0.284000 0.298000 0.376000 0.733000 ;
        RECT 0.049000 0.652000 0.376000 0.733000 ;
        RECT 0.049000 0.298000 0.376000 0.379000 ;
    END
END BUFX4

MACRO BUFX3
    CLASS CORE ;
    FOREIGN BUFX3 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 0.700000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.037000 0.433000 0.147000 0.562000 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 0.700000 1.280000 ;
        RECT 0.196000 1.078000 0.286000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 0.700000 0.080000 ;
        RECT 0.557000 -0.080000 0.647000 0.122000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.387000 0.433000 0.488000 0.633000 ;
        RECT 0.398000 0.433000 0.488000 0.752000 ;
        RECT 0.408000 0.287000 0.498000 0.368000 ;
        RECT 0.408000 0.287000 0.469000 0.752000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 0.235000 0.470000 0.325000 0.551000 ;
        RECT 0.048000 0.696000 0.138000 0.777000 ;
        RECT 0.048000 0.244000 0.138000 0.325000 ;
        RECT 0.235000 0.270000 0.296000 0.751000 ;
        RECT 0.048000 0.696000 0.296000 0.751000 ;
        RECT 0.048000 0.270000 0.296000 0.325000 ;
    END
END BUFX3

MACRO BUFX2
    CLASS CORE ;
    FOREIGN BUFX2 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 0.700000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.037000 0.418000 0.236000 0.538000 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 0.700000 1.280000 ;
        RECT 0.223000 1.078000 0.313000 1.280000 ;
        RECT 0.237000 1.065000 0.298000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 0.700000 0.080000 ;
        RECT 0.233000 -0.080000 0.323000 0.122000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.435000 0.331000 0.525000 0.412000 ;
        RECT 0.424000 0.655000 0.514000 0.736000 ;
        RECT 0.562000 0.357000 0.623000 0.710000 ;
        RECT 0.562000 0.439000 0.643000 0.494000 ;
        RECT 0.435000 0.357000 0.623000 0.412000 ;
        RECT 0.424000 0.655000 0.623000 0.710000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 0.302000 0.490000 0.430000 0.571000 ;
        RECT 0.074000 0.657000 0.164000 0.738000 ;
        RECT 0.074000 0.275000 0.164000 0.356000 ;
        RECT 0.302000 0.301000 0.363000 0.712000 ;
        RECT 0.074000 0.657000 0.363000 0.712000 ;
        RECT 0.074000 0.301000 0.363000 0.356000 ;
    END
END BUFX2

MACRO BUFX12
    CLASS CORE ;
    FOREIGN BUFX12 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 1.800000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.194000 0.474000 0.554000 0.555000 ;
        RECT 0.239000 0.439000 0.301000 0.555000 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 1.800000 1.280000 ;
        RECT 1.658000 0.972000 1.751000 1.280000 ;
        RECT 0.922000 0.972000 1.015000 1.280000 ;
        RECT 1.285000 0.972000 1.377000 1.280000 ;
        RECT 0.573000 0.897000 0.665000 1.280000 ;
        RECT 0.224000 0.897000 0.316000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 1.800000 0.080000 ;
        RECT 1.642000 -0.080000 1.735000 0.211000 ;
        RECT 1.293000 -0.080000 1.385000 0.211000 ;
        RECT 0.944000 -0.080000 1.036000 0.215000 ;
        RECT 0.595000 -0.080000 0.687000 0.215000 ;
        RECT 0.235000 -0.080000 0.327000 0.122000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.319000 0.300000 1.741000 0.767000 ;
        RECT 1.298000 0.626000 1.741000 0.757000 ;
        RECT 1.298000 0.321000 1.741000 0.440000 ;
        RECT 0.769000 0.321000 1.741000 0.402000 ;
        RECT 0.747000 0.676000 1.741000 0.757000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 0.622000 0.519000 1.193000 0.600000 ;
        RECT 0.420000 0.319000 0.513000 0.400000 ;
        RECT 0.398000 0.657000 0.491000 0.738000 ;
        RECT 0.049000 0.657000 0.142000 0.738000 ;
        RECT 0.622000 0.345000 0.685000 0.712000 ;
        RECT 0.079000 0.319000 0.142000 0.389000 ;
        RECT 0.420000 0.345000 0.685000 0.400000 ;
        RECT 0.079000 0.319000 0.513000 0.374000 ;
        RECT 0.049000 0.657000 0.685000 0.712000 ;
        RECT 0.049000 0.335000 0.142000 0.389000 ;
    END
END BUFX12

MACRO AOI33X2
    CLASS CORE ;
    FOREIGN AOI33X2 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 2.300000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.541000 0.525000 1.732000 0.633000 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.351000 0.411000 1.413000 0.640000 ;
        RECT 1.815000 0.411000 1.876000 0.574000 ;
        RECT 1.351000 0.411000 1.876000 0.465000 ;
        RECT 1.296000 0.573000 1.413000 0.627000 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 2.037000 0.301000 2.099000 0.481000 ;
        RECT 1.137000 0.301000 1.198000 0.554000 ;
        RECT 1.137000 0.301000 2.099000 0.356000 ;
        RECT 1.119000 0.439000 1.198000 0.494000 ;
        END
    END A2
    PIN B0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.477000 0.439000 0.578000 0.540000 ;
        RECT 0.411000 0.439000 0.578000 0.494000 ;
        END
    END B0
    PIN B1
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.765000 0.439000 0.827000 0.650000 ;
        RECT 0.294000 0.595000 0.878000 0.650000 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.969000 0.679000 1.071000 0.760000 ;
        RECT 0.126000 0.573000 0.188000 0.760000 ;
        RECT 0.126000 0.705000 1.071000 0.760000 ;
        RECT 0.058000 0.573000 0.188000 0.627000 ;
        END
    END B2
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 2.300000 1.280000 ;
        RECT 0.906000 0.984000 0.997000 1.280000 ;
        RECT 0.563000 0.984000 0.654000 1.280000 ;
        RECT 0.220000 0.984000 0.311000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 2.300000 0.080000 ;
        RECT 2.055000 -0.080000 2.146000 0.122000 ;
        RECT 1.047000 -0.080000 1.138000 0.122000 ;
        RECT 0.048000 -0.080000 0.139000 0.403000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 2.161000 0.192000 2.242000 0.306000 ;
        RECT 2.181000 0.192000 2.242000 0.787000 ;
        RECT 0.885000 0.192000 0.946000 0.352000 ;
        RECT 1.272000 0.732000 2.242000 0.787000 ;
        RECT 0.885000 0.192000 2.242000 0.246000 ;
        RECT 0.541000 0.298000 0.946000 0.352000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 2.132000 0.896000 2.224000 0.977000 ;
        RECT 1.787000 0.896000 1.878000 0.977000 ;
        RECT 1.444000 0.896000 1.535000 0.977000 ;
        RECT 1.100000 0.896000 1.192000 0.977000 ;
        RECT 1.100000 0.814000 1.162000 0.977000 ;
        RECT 0.048000 0.814000 1.162000 0.869000 ;
        RECT 1.878000 0.910000 2.132000 0.964000 ;
        RECT 1.535000 0.910000 1.787000 0.964000 ;
        RECT 1.192000 0.910000 1.444000 0.964000 ;
    END
END AOI33X2

MACRO AOI32X2
    CLASS CORE ;
    FOREIGN AOI32X2 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 2.000000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.490000 0.306000 0.554000 0.468000 ;
        RECT 0.490000 0.413000 0.584000 0.468000 ;
        RECT 0.423000 0.306000 0.554000 0.361000 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.766000 0.439000 0.872000 0.577000 ;
        RECT 0.302000 0.523000 0.872000 0.577000 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.948000 0.626000 1.056000 0.692000 ;
        RECT 0.114000 0.573000 0.178000 0.692000 ;
        RECT 0.993000 0.569000 1.056000 0.692000 ;
        RECT 0.114000 0.637000 1.056000 0.692000 ;
        RECT 0.059000 0.573000 0.178000 0.627000 ;
        END
    END A2
    PIN B0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.372000 0.433000 1.466000 0.550000 ;
        RECT 1.371000 0.433000 1.598000 0.507000 ;
        END
    END B0
    PIN B1
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.150000 0.439000 1.241000 0.507000 ;
        RECT 1.178000 0.439000 1.241000 0.661000 ;
        RECT 1.178000 0.606000 1.742000 0.661000 ;
        END
    END B1
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 2.000000 1.280000 ;
        RECT 0.580000 0.989000 0.674000 1.280000 ;
        RECT 0.226000 0.989000 0.320000 1.280000 ;
        RECT 0.933000 0.989000 1.026000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 2.000000 0.080000 ;
        RECT 1.074000 -0.080000 1.168000 0.122000 ;
        RECT 1.791000 -0.080000 1.884000 0.275000 ;
        RECT 0.065000 -0.080000 0.128000 0.325000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.857000 0.348000 1.941000 0.439000 ;
        RECT 1.663000 0.721000 1.756000 0.802000 ;
        RECT 1.310000 0.719000 1.404000 0.800000 ;
        RECT 1.877000 0.348000 1.941000 0.789000 ;
        RECT 1.664000 0.281000 1.727000 0.402000 ;
        RECT 0.831000 0.189000 0.894000 0.336000 ;
        RECT 1.310000 0.732000 1.756000 0.787000 ;
        RECT 0.831000 0.281000 1.727000 0.336000 ;
        RECT 0.556000 0.189000 0.894000 0.244000 ;
        RECT 1.664000 0.348000 1.941000 0.402000 ;
        RECT 1.663000 0.735000 1.941000 0.789000 ;
        RECT 1.310000 0.735000 1.941000 0.787000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 1.839000 0.896000 1.933000 0.977000 ;
        RECT 1.486000 0.896000 1.580000 0.977000 ;
        RECT 1.134000 0.896000 1.227000 0.977000 ;
        RECT 0.756000 0.799000 0.850000 0.880000 ;
        RECT 0.404000 0.796000 0.497000 0.877000 ;
        RECT 0.050000 0.796000 0.143000 0.877000 ;
        RECT 1.134000 0.812000 1.197000 0.977000 ;
        RECT 0.850000 0.812000 1.134000 0.867000 ;
        RECT 1.580000 0.910000 1.839000 0.964000 ;
        RECT 1.227000 0.910000 1.486000 0.964000 ;
        RECT 0.497000 0.810000 0.756000 0.864000 ;
        RECT 0.143000 0.810000 0.404000 0.864000 ;
    END
END AOI32X2

MACRO AOI31X4
    CLASS CORE ;
    FOREIGN AOI31X4 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 1.600000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.381000 0.410000 0.521000 0.507000 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.201000 0.567000 0.341000 0.726000 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.038000 0.363000 0.140000 0.500000 ;
        END
    END A2
    PIN B0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.707000 0.429000 0.851000 0.564000 ;
        END
    END B0
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 1.600000 1.280000 ;
        RECT 0.350000 1.078000 0.442000 1.280000 ;
        RECT 0.048000 1.078000 0.140000 1.280000 ;
        RECT 1.090000 0.910000 1.181000 1.280000 ;
        RECT 1.451000 0.904000 1.512000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 1.600000 0.080000 ;
        RECT 0.048000 -0.080000 0.140000 0.292000 ;
        RECT 1.436000 -0.080000 1.527000 0.214000 ;
        RECT 1.090000 -0.080000 1.181000 0.214000 ;
        RECT 0.706000 -0.080000 0.797000 0.122000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.460000 0.433000 1.562000 0.767000 ;
        RECT 1.460000 0.337000 1.546000 0.767000 ;
        RECT 1.262000 0.337000 1.546000 0.392000 ;
        RECT 1.263000 0.667000 1.562000 0.721000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 1.040000 0.485000 1.397000 0.571000 ;
        RECT 0.559000 0.265000 0.645000 0.354000 ;
        RECT 1.040000 0.313000 1.102000 0.818000 ;
        RECT 0.929000 0.763000 0.991000 1.042000 ;
        RECT 0.913000 0.443000 0.975000 0.698000 ;
        RECT 0.909000 0.152000 0.971000 0.368000 ;
        RECT 0.764000 0.643000 0.826000 0.867000 ;
        RECT 0.583000 0.265000 0.645000 0.698000 ;
        RECT 0.929000 0.763000 1.102000 0.818000 ;
        RECT 0.909000 0.313000 1.102000 0.368000 ;
        RECT 0.896000 0.987000 0.991000 1.042000 ;
        RECT 0.583000 0.643000 0.975000 0.698000 ;
        RECT 0.199000 0.839000 0.646000 0.894000 ;
    END
END AOI31X4

MACRO AOI31X2
    CLASS CORE ;
    FOREIGN AOI31X2 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 1.600000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.038000 0.550000 0.140000 0.692000 ;
        RECT 0.990000 0.490000 1.052000 0.692000 ;
        RECT 0.038000 0.637000 1.052000 0.692000 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.749000 0.439000 0.851000 0.582000 ;
        RECT 0.329000 0.527000 0.882000 0.582000 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.236000 0.306000 0.318000 0.468000 ;
        RECT 0.236000 0.413000 0.614000 0.468000 ;
        END
    END A2
    PIN B0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.248000 0.433000 1.395000 0.557000 ;
        END
    END B0
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 1.600000 1.280000 ;
        RECT 0.910000 0.911000 1.002000 1.280000 ;
        RECT 0.566000 0.911000 0.657000 1.280000 ;
        RECT 0.221000 0.911000 0.312000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 1.600000 0.080000 ;
        RECT 1.244000 -0.080000 1.336000 0.122000 ;
        RECT 0.544000 -0.080000 0.636000 0.198000 ;
        RECT 1.269000 -0.080000 1.331000 0.304000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.282000 0.627000 1.354000 0.706000 ;
        RECT 1.292000 0.627000 1.354000 0.800000 ;
        RECT 1.125000 0.268000 1.187000 0.682000 ;
        RECT 0.420000 0.158000 0.482000 0.323000 ;
        RECT 1.125000 0.627000 1.354000 0.682000 ;
        RECT 0.420000 0.268000 1.187000 0.323000 ;
        RECT 0.048000 0.158000 0.482000 0.213000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 1.067000 0.746000 1.129000 0.964000 ;
        RECT 0.048000 0.746000 1.129000 0.801000 ;
        RECT 1.067000 0.910000 1.541000 0.964000 ;
    END
END AOI31X2

MACRO AOI2BB2X2
    CLASS CORE ;
    FOREIGN AOI2BB2X2 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 1.600000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A0N
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.038000 0.445000 0.140000 0.633000 ;
        END
    END A0N
    PIN A1N
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.343000 0.388000 0.496000 0.500000 ;
        END
    END A1N
    PIN B0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.294000 0.379000 1.371000 0.498000 ;
        RECT 0.672000 0.379000 1.371000 0.433000 ;
        END
    END B0
    PIN B1
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.104000 0.543000 1.201000 0.737000 ;
        RECT 0.512000 0.682000 1.201000 0.737000 ;
        END
    END B1
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 1.600000 1.280000 ;
        RECT 1.449000 1.078000 1.541000 1.280000 ;
        RECT 0.404000 0.988000 0.496000 1.280000 ;
        RECT 0.749000 0.988000 0.840000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 1.600000 0.080000 ;
        RECT 0.980000 -0.080000 1.072000 0.122000 ;
        RECT 0.424000 -0.080000 0.516000 0.289000 ;
        RECT 0.048000 -0.080000 0.140000 0.122000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.203000 0.923000 1.304000 1.040000 ;
        RECT 1.187000 0.967000 1.304000 1.040000 ;
        RECT 1.446000 0.192000 1.508000 0.977000 ;
        RECT 1.446000 0.306000 1.542000 0.361000 ;
        RECT 1.203000 0.923000 1.508000 0.977000 ;
        RECT 1.094000 0.986000 1.304000 1.040000 ;
        RECT 0.773000 0.192000 1.508000 0.246000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 0.214000 0.288000 0.276000 0.788000 ;
        RECT 0.576000 0.808000 1.358000 0.863000 ;
        RECT 0.214000 0.571000 0.991000 0.626000 ;
        RECT 0.048000 0.733000 0.276000 0.788000 ;
    END
END AOI2BB2X2

MACRO AOI2BB1X4
    CLASS CORE ;
    FOREIGN AOI2BB1X4 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 2.000000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A0N
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.271000 0.439000 0.335000 0.648000 ;
        RECT 0.241000 0.439000 0.335000 0.494000 ;
        END
    END A0N
    PIN A1N
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.067000 0.567000 0.131000 0.889000 ;
        RECT 0.594000 0.439000 0.657000 0.889000 ;
        RECT 0.594000 0.439000 0.668000 0.494000 ;
        RECT 0.067000 0.835000 0.657000 0.889000 ;
        END
    END A1N
    PIN B0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.785000 0.433000 0.893000 0.602000 ;
        END
    END B0
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 2.000000 1.280000 ;
        RECT 0.667000 1.078000 0.760000 1.280000 ;
        RECT 0.050000 1.078000 0.143000 1.280000 ;
        RECT 1.365000 0.973000 1.428000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 2.000000 0.080000 ;
        RECT 1.702000 -0.080000 1.796000 0.122000 ;
        RECT 1.267000 -0.080000 1.361000 0.198000 ;
        RECT 0.861000 -0.080000 0.955000 0.198000 ;
        RECT 0.468000 -0.080000 0.562000 0.198000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.493000 0.700000 1.618000 0.894000 ;
        RECT 1.493000 0.700000 1.598000 1.033000 ;
        RECT 1.493000 0.700000 1.697000 0.767000 ;
        RECT 1.555000 0.318000 1.618000 0.894000 ;
        RECT 1.084000 0.318000 1.147000 0.412000 ;
        RECT 1.084000 0.318000 1.618000 0.373000 ;
        RECT 1.019000 0.706000 1.774000 0.761000 ;
        RECT 1.555000 0.318000 1.598000 1.033000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 1.428000 0.458000 1.492000 0.630000 ;
        RECT 0.956000 0.324000 1.019000 0.630000 ;
        RECT 0.398000 0.324000 0.461000 0.761000 ;
        RECT 0.956000 0.575000 1.492000 0.630000 ;
        RECT 0.358000 0.706000 0.461000 0.761000 ;
        RECT 0.269000 0.324000 1.019000 0.379000 ;
    END
END AOI2BB1X4

MACRO AOI2BB1X2
    CLASS CORE ;
    FOREIGN AOI2BB1X2 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 1.300000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A0N
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.039000 0.300000 0.149000 0.429000 ;
        END
    END A0N
    PIN A1N
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.194000 0.555000 0.387000 0.652000 ;
        END
    END A1N
    PIN B0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.606000 0.439000 0.671000 0.538000 ;
        RECT 1.009000 0.439000 1.073000 0.638000 ;
        RECT 0.606000 0.439000 1.073000 0.494000 ;
        END
    END B0
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 1.300000 1.280000 ;
        RECT 1.097000 0.860000 1.193000 1.280000 ;
        RECT 0.366000 1.078000 0.461000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 1.300000 0.080000 ;
        RECT 0.872000 -0.080000 0.968000 0.122000 ;
        RECT 0.456000 -0.080000 0.552000 0.198000 ;
        RECT 0.051000 -0.080000 0.146000 0.198000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.737000 0.711000 0.868000 0.894000 ;
        RECT 0.737000 0.711000 0.833000 0.904000 ;
        RECT 0.674000 0.300000 0.803000 0.377000 ;
        RECT 0.674000 0.162000 0.739000 0.377000 ;
        RECT 1.147000 0.323000 1.211000 0.765000 ;
        RECT 0.737000 0.711000 1.211000 0.765000 ;
        RECT 0.674000 0.323000 1.211000 0.377000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 0.051000 0.707000 0.146000 0.900000 ;
        RECT 0.453000 0.427000 0.518000 0.762000 ;
        RECT 0.269000 0.183000 0.333000 0.482000 ;
        RECT 0.453000 0.596000 0.900000 0.651000 ;
        RECT 0.269000 0.427000 0.518000 0.482000 ;
        RECT 0.051000 0.707000 0.518000 0.762000 ;
    END
END AOI2BB1X2

MACRO AOI22X2
    CLASS CORE ;
    FOREIGN AOI22X2 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 1.600000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.061000 0.567000 1.207000 0.661000 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.356000 0.438000 1.418000 0.551000 ;
        RECT 0.882000 0.438000 0.944000 0.664000 ;
        RECT 0.882000 0.438000 1.009000 0.494000 ;
        RECT 0.882000 0.438000 1.418000 0.493000 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.329000 0.573000 0.475000 0.663000 ;
        END
    END B0
    PIN B1
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.185000 0.439000 0.298000 0.511000 ;
        RECT 0.113000 0.493000 0.246000 0.562000 ;
        RECT 0.653000 0.456000 0.715000 0.575000 ;
        RECT 0.185000 0.439000 0.246000 0.562000 ;
        RECT 0.185000 0.456000 0.715000 0.511000 ;
        END
    END B1
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 1.600000 1.280000 ;
        RECT 0.566000 0.888000 0.657000 1.280000 ;
        RECT 0.221000 0.888000 0.312000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 1.600000 0.080000 ;
        RECT 1.352000 -0.080000 1.444000 0.122000 ;
        RECT 0.695000 -0.080000 0.787000 0.122000 ;
        RECT 0.048000 -0.080000 0.140000 0.305000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.302000 0.706000 1.368000 0.789000 ;
        RECT 1.480000 0.321000 1.542000 0.761000 ;
        RECT 1.302000 0.706000 1.542000 0.761000 ;
        RECT 0.393000 0.321000 1.542000 0.376000 ;
        RECT 0.932000 0.735000 1.368000 0.789000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 0.753000 0.732000 0.815000 0.940000 ;
        RECT 0.048000 0.732000 0.830000 0.787000 ;
        RECT 0.753000 0.886000 1.541000 0.940000 ;
    END
END AOI22X2

MACRO AOI222X4
    CLASS CORE ;
    FOREIGN AOI222X4 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 2.100000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.912000 0.398000 1.013000 0.556000 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.094000 0.524000 1.188000 0.686000 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.737000 0.505000 0.838000 0.777000 ;
        END
    END B0
    PIN B1
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.407000 0.573000 0.642000 0.627000 ;
        END
    END B1
    PIN C0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.231000 0.382000 0.414000 0.494000 ;
        END
    END C0
    PIN C1
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.037000 0.433000 0.138000 0.624000 ;
        END
    END C1
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 2.100000 1.280000 ;
        RECT 1.893000 0.982000 1.983000 1.280000 ;
        RECT 1.554000 0.908000 1.644000 1.280000 ;
        RECT 0.345000 1.078000 0.435000 1.280000 ;
        RECT 0.048000 1.078000 0.138000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 2.100000 0.080000 ;
        RECT 0.048000 -0.080000 0.180000 0.083000 ;
        RECT 1.893000 -0.080000 1.983000 0.212000 ;
        RECT 1.543000 -0.080000 1.633000 0.212000 ;
        RECT 1.167000 -0.080000 1.257000 0.122000 ;
        RECT 0.573000 -0.080000 0.663000 0.122000 ;
        RECT 0.048000 -0.080000 0.138000 0.275000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.787000 0.567000 1.888000 0.900000 ;
        RECT 1.787000 0.336000 1.875000 0.440000 ;
        RECT 1.723000 0.661000 1.888000 0.742000 ;
        RECT 1.814000 0.336000 1.875000 0.900000 ;
        RECT 1.723000 0.336000 1.875000 0.390000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 0.870000 0.236000 0.963000 0.320000 ;
        RECT 1.534000 0.287000 1.595000 0.705000 ;
        RECT 1.377000 0.650000 1.438000 0.740000 ;
        RECT 1.249000 0.404000 1.310000 0.833000 ;
        RECT 1.078000 0.265000 1.139000 0.458000 ;
        RECT 1.534000 0.530000 1.725000 0.585000 ;
        RECT 1.377000 0.650000 1.595000 0.705000 ;
        RECT 1.352000 0.287000 1.595000 0.342000 ;
        RECT 1.249000 0.520000 1.450000 0.575000 ;
        RECT 0.870000 0.265000 1.139000 0.320000 ;
        RECT 0.530000 0.995000 1.267000 1.050000 ;
        RECT 0.196000 0.812000 0.639000 0.867000 ;
        RECT 1.078000 0.404000 1.310000 0.458000 ;
        RECT 1.029000 0.779000 1.310000 0.833000 ;
        RECT 0.387000 0.236000 0.963000 0.290000 ;
    END
END AOI222X4

MACRO AOI222X2
    CLASS CORE ;
    FOREIGN AOI222X2 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 2.500000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.814000 0.556000 2.016000 0.627000 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 2.210000 0.439000 2.273000 0.545000 ;
        RECT 1.665000 0.439000 2.273000 0.494000 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.130000 0.558000 1.331000 0.627000 ;
        END
    END B0
    PIN B1
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.951000 0.439000 1.558000 0.494000 ;
        END
    END B1
    PIN C0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.319000 0.398000 0.517000 0.507000 ;
        END
    END C0
    PIN C1
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.628000 0.556000 0.725000 0.620000 ;
        RECT 0.093000 0.521000 0.156000 0.627000 ;
        RECT 0.093000 0.565000 0.299000 0.627000 ;
        RECT 0.093000 0.565000 0.725000 0.620000 ;
        END
    END C1
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 2.500000 1.280000 ;
        RECT 0.741000 0.911000 0.833000 1.280000 ;
        RECT 0.395000 0.911000 0.487000 1.280000 ;
        RECT 0.049000 0.911000 0.141000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 2.500000 0.080000 ;
        RECT 2.261000 -0.080000 2.353000 0.198000 ;
        RECT 1.567000 -0.080000 1.659000 0.198000 ;
        RECT 0.782000 -0.080000 0.874000 0.198000 ;
        RECT 0.049000 -0.080000 0.141000 0.275000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 2.263000 0.268000 2.399000 0.367000 ;
        RECT 1.905000 0.249000 2.024000 0.323000 ;
        RECT 1.190000 0.249000 1.318000 0.323000 ;
        RECT 2.336000 0.268000 2.399000 0.743000 ;
        RECT 2.201000 0.688000 2.263000 0.761000 ;
        RECT 1.797000 0.688000 2.399000 0.743000 ;
        RECT 0.395000 0.268000 2.399000 0.323000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 0.222000 0.688000 1.542000 0.743000 ;
        RECT 0.931000 0.910000 2.408000 0.964000 ;
    END
END AOI222X2

MACRO AOI221X4
    CLASS CORE ;
    FOREIGN AOI221X4 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 2.000000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.423000 0.433000 0.534000 0.585000 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.668000 0.502000 0.731000 0.627000 ;
        RECT 0.668000 0.567000 0.850000 0.627000 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.241000 0.598000 0.336000 0.761000 ;
        END
    END B0
    PIN B1
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.039000 0.462000 0.143000 0.632000 ;
        END
    END B1
    PIN C0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.862000 0.373000 1.032000 0.494000 ;
        END
    END C0
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 2.000000 1.280000 ;
        RECT 1.840000 0.765000 1.934000 1.280000 ;
        RECT 0.358000 1.078000 0.452000 1.280000 ;
        RECT 1.444000 0.765000 1.537000 1.280000 ;
        RECT 0.050000 1.078000 0.143000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 2.000000 0.080000 ;
        RECT 1.427000 -0.080000 1.521000 0.198000 ;
        RECT 0.766000 -0.080000 0.860000 0.122000 ;
        RECT 0.050000 -0.080000 0.143000 0.291000 ;
        RECT 1.843000 -0.080000 1.906000 0.361000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.675000 0.300000 1.780000 0.633000 ;
        RECT 1.642000 0.660000 1.738000 0.964000 ;
        RECT 1.675000 0.300000 1.738000 0.964000 ;
        RECT 1.625000 0.300000 1.780000 0.355000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 1.084000 0.723000 1.179000 0.810000 ;
        RECT 1.245000 0.895000 1.339000 0.976000 ;
        RECT 1.333000 0.345000 1.397000 0.644000 ;
        RECT 1.275000 0.589000 1.339000 0.976000 ;
        RECT 1.242000 0.274000 1.306000 0.400000 ;
        RECT 1.116000 0.236000 1.179000 0.810000 ;
        RECT 0.602000 0.236000 0.665000 0.306000 ;
        RECT 1.333000 0.508000 1.573000 0.563000 ;
        RECT 1.275000 0.589000 1.397000 0.644000 ;
        RECT 1.242000 0.345000 1.397000 0.400000 ;
        RECT 1.116000 0.468000 1.270000 0.523000 ;
        RECT 0.402000 0.251000 0.665000 0.306000 ;
        RECT 0.204000 0.832000 0.799000 0.887000 ;
        RECT 0.602000 0.236000 1.179000 0.290000 ;
        RECT 1.333000 0.345000 1.339000 0.976000 ;
    END
END AOI221X4

MACRO AOI221X2
    CLASS CORE ;
    FOREIGN AOI221X2 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 2.100000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.087000 0.396000 1.233000 0.500000 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.932000 0.573000 0.993000 0.650000 ;
        RECT 0.917000 0.595000 1.572000 0.650000 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.212000 0.306000 0.313000 0.430000 ;
        RECT 0.212000 0.375000 0.414000 0.430000 ;
        END
    END B0
    PIN B1
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.562000 0.433000 0.663000 0.558000 ;
        RECT 0.562000 0.493000 0.711000 0.558000 ;
        RECT 0.077000 0.504000 0.711000 0.558000 ;
        END
    END B1
    PIN C0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.678000 0.439000 1.739000 0.543000 ;
        RECT 1.457000 0.439000 1.739000 0.494000 ;
        END
    END C0
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 2.100000 1.280000 ;
        RECT 0.727000 0.903000 0.817000 1.280000 ;
        RECT 0.387000 0.903000 0.477000 1.280000 ;
        RECT 0.048000 0.903000 0.138000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 2.100000 0.080000 ;
        RECT 1.546000 -0.080000 1.636000 0.198000 ;
        RECT 0.780000 -0.080000 0.870000 0.122000 ;
        RECT 0.048000 -0.080000 0.138000 0.198000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.761000 0.755000 1.868000 0.836000 ;
        RECT 1.330000 0.300000 1.457000 0.367000 ;
        RECT 1.807000 0.312000 1.868000 0.836000 ;
        RECT 1.330000 0.225000 1.391000 0.367000 ;
        RECT 1.330000 0.312000 1.868000 0.367000 ;
        RECT 0.387000 0.225000 1.391000 0.280000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 0.883000 0.707000 0.944000 0.823000 ;
        RECT 0.912000 0.962000 2.020000 1.017000 ;
        RECT 0.883000 0.768000 1.511000 0.823000 ;
        RECT 0.217000 0.707000 0.944000 0.762000 ;
    END
END AOI221X2

MACRO AOI21X4
    CLASS CORE ;
    FOREIGN AOI21X4 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 1.800000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.115000 0.469000 0.207000 0.574000 ;
        RECT 0.745000 0.530000 0.807000 0.627000 ;
        RECT 0.145000 0.469000 0.207000 0.625000 ;
        RECT 0.145000 0.567000 0.218000 0.625000 ;
        RECT 0.145000 0.570000 0.807000 0.625000 ;
        RECT 0.745000 0.573000 0.841000 0.627000 ;
        RECT 0.145000 0.573000 0.841000 0.625000 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.415000 0.392000 0.661000 0.494000 ;
        RECT 1.005000 0.452000 1.098000 0.533000 ;
        RECT 0.400000 0.426000 0.492000 0.507000 ;
        RECT 0.415000 0.392000 0.492000 0.507000 ;
        RECT 0.400000 0.426000 0.661000 0.494000 ;
        RECT 1.005000 0.392000 1.068000 0.533000 ;
        RECT 0.415000 0.392000 1.068000 0.446000 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.238000 0.496000 1.402000 0.635000 ;
        END
    END B0
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 1.800000 1.280000 ;
        RECT 0.922000 0.941000 1.015000 1.280000 ;
        RECT 0.573000 0.941000 0.665000 1.280000 ;
        RECT 0.224000 0.941000 0.316000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 1.800000 0.080000 ;
        RECT 1.458000 -0.080000 1.550000 0.122000 ;
        RECT 1.098000 -0.080000 1.190000 0.198000 ;
        RECT 0.400000 -0.080000 0.492000 0.198000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.208000 0.274000 1.319000 0.392000 ;
        RECT 1.478000 0.300000 1.582000 0.633000 ;
        RECT 1.620000 0.896000 1.713000 0.977000 ;
        RECT 1.271000 0.896000 1.364000 0.977000 ;
        RECT 1.605000 0.896000 1.713000 0.964000 ;
        RECT 1.605000 0.579000 1.668000 0.964000 ;
        RECT 1.208000 0.337000 1.582000 0.392000 ;
        RECT 0.049000 0.274000 1.319000 0.329000 ;
        RECT 1.478000 0.579000 1.668000 0.633000 ;
        RECT 1.271000 0.910000 1.713000 0.964000 ;
        RECT 1.620000 0.579000 1.668000 0.977000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 0.049000 0.698000 1.538000 0.752000 ;
    END
END AOI21X4

MACRO AOI21X2
    CLASS CORE ;
    FOREIGN AOI21X2 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 1.300000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.039000 0.433000 0.146000 0.530000 ;
        RECT 0.039000 0.457000 0.763000 0.512000 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.246000 0.595000 0.518000 0.669000 ;
        RECT 0.246000 0.573000 0.311000 0.669000 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.830000 0.485000 0.936000 0.627000 ;
        RECT 0.803000 0.573000 0.936000 0.627000 ;
        END
    END B0
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 1.300000 1.280000 ;
        RECT 0.591000 0.888000 0.687000 1.280000 ;
        RECT 0.231000 0.888000 0.326000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 1.300000 0.080000 ;
        RECT 0.986000 -0.080000 1.082000 0.122000 ;
        RECT 0.411000 -0.080000 0.506000 0.275000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.771000 0.268000 0.867000 0.400000 ;
        RECT 0.989000 0.706000 1.095000 0.789000 ;
        RECT 0.051000 0.268000 0.146000 0.349000 ;
        RECT 1.030000 0.345000 1.095000 0.789000 ;
        RECT 0.235000 0.294000 0.300000 0.400000 ;
        RECT 0.235000 0.345000 1.095000 0.400000 ;
        RECT 0.051000 0.294000 0.300000 0.349000 ;
        RECT 0.974000 0.735000 1.095000 0.789000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 1.154000 0.873000 1.249000 0.954000 ;
        RECT 0.806000 0.732000 0.871000 0.927000 ;
        RECT 0.051000 0.732000 0.871000 0.787000 ;
        RECT 0.806000 0.873000 1.249000 0.927000 ;
    END
END AOI21X2

MACRO AND4X4
    CLASS CORE ;
    FOREIGN AND4X4 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 2.000000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.579000 0.625000 0.689000 0.773000 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.766000 0.489000 0.871000 0.629000 ;
        RECT 0.460000 0.489000 0.871000 0.544000 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.220000 0.493000 0.344000 0.636000 ;
        RECT 0.220000 0.539000 0.364000 0.636000 ;
        RECT 0.988000 0.379000 1.051000 0.721000 ;
        RECT 0.281000 0.379000 0.344000 0.636000 ;
        RECT 0.948000 0.379000 1.051000 0.439000 ;
        RECT 0.281000 0.379000 1.051000 0.433000 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.039000 0.640000 0.146000 0.767000 ;
        RECT 1.213000 0.567000 1.328000 0.650000 ;
        RECT 1.264000 0.439000 1.328000 0.650000 ;
        RECT 1.114000 0.595000 1.178000 0.888000 ;
        RECT 0.081000 0.640000 0.145000 0.888000 ;
        RECT 1.264000 0.439000 1.364000 0.494000 ;
        RECT 1.114000 0.595000 1.328000 0.650000 ;
        RECT 0.081000 0.833000 1.178000 0.888000 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 2.000000 1.280000 ;
        RECT 1.643000 1.078000 1.751000 1.280000 ;
        RECT 0.251000 1.078000 0.358000 1.280000 ;
        RECT 1.131000 1.078000 1.225000 1.280000 ;
        RECT 0.689000 1.078000 0.782000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 2.000000 0.080000 ;
        RECT 1.372000 -0.080000 1.466000 0.250000 ;
        RECT 1.769000 -0.080000 1.862000 0.211000 ;
        RECT 0.050000 -0.080000 0.143000 0.334000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.675000 0.567000 1.780000 0.900000 ;
        RECT 1.438000 0.815000 1.532000 1.039000 ;
        RECT 1.438000 0.815000 1.780000 0.900000 ;
        RECT 1.676000 0.356000 1.759000 0.900000 ;
        RECT 1.675000 0.356000 1.759000 0.439000 ;
        RECT 1.570000 0.331000 1.696000 0.412000 ;
        RECT 1.570000 0.356000 1.759000 0.412000 ;
        RECT 1.676000 0.331000 1.696000 0.900000 ;
        RECT 1.675000 0.331000 1.676000 0.439000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 0.905000 0.944000 0.999000 1.039000 ;
        RECT 0.479000 0.944000 0.573000 1.039000 ;
        RECT 1.444000 0.507000 1.574000 0.588000 ;
        RECT 0.711000 0.240000 0.804000 0.321000 ;
        RECT 1.242000 0.706000 1.306000 0.999000 ;
        RECT 1.444000 0.329000 1.507000 0.761000 ;
        RECT 1.164000 0.254000 1.227000 0.383000 ;
        RECT 1.242000 0.706000 1.507000 0.761000 ;
        RECT 0.479000 0.944000 1.306000 0.999000 ;
        RECT 1.164000 0.329000 1.507000 0.383000 ;
        RECT 0.905000 0.254000 1.227000 0.308000 ;
        RECT 0.804000 0.254000 1.164000 0.308000 ;
        RECT 0.711000 0.254000 0.999000 0.308000 ;
    END
END AND4X4

MACRO AND4X2
    CLASS CORE ;
    FOREIGN AND4X2 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 1.100000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.039000 0.398000 0.157000 0.556000 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.222000 0.537000 0.358000 0.645000 ;
        RECT 0.279000 0.537000 0.358000 0.646000 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.478000 0.581000 0.542000 0.761000 ;
        RECT 0.426000 0.706000 0.542000 0.761000 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.610000 0.439000 0.694000 0.606000 ;
        RECT 0.610000 0.524000 0.733000 0.606000 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 1.100000 1.280000 ;
        RECT 0.724000 1.064000 0.838000 1.280000 ;
        RECT 0.049000 1.078000 0.158000 1.280000 ;
        RECT 0.419000 1.078000 0.514000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 1.100000 0.080000 ;
        RECT 0.721000 -0.080000 0.815000 0.122000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.967000 0.648000 1.049000 0.767000 ;
        RECT 0.967000 0.700000 1.061000 0.767000 ;
        RECT 0.985000 0.358000 1.049000 0.767000 ;
        RECT 0.967000 0.648000 1.031000 0.964000 ;
        RECT 0.967000 0.199000 1.031000 0.413000 ;
        RECT 0.967000 0.358000 1.049000 0.413000 ;
        RECT 0.985000 0.199000 1.031000 0.964000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 0.061000 0.250000 0.156000 0.343000 ;
        RECT 0.825000 0.473000 0.919000 0.556000 ;
        RECT 0.076000 0.211000 0.156000 0.343000 ;
        RECT 0.825000 0.211000 0.889000 0.889000 ;
        RECT 0.208000 0.835000 0.889000 0.889000 ;
        RECT 0.076000 0.211000 0.889000 0.265000 ;
    END
END AND4X2

MACRO AOI211X2
    CLASS CORE ;
    FOREIGN AOI211X2 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 1.600000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.524000 0.540000 0.615000 0.621000 ;
        RECT 0.116000 0.386000 0.207000 0.467000 ;
        RECT 0.539000 0.494000 0.615000 0.621000 ;
        RECT 0.058000 0.399000 0.207000 0.467000 ;
        RECT 0.539000 0.399000 0.601000 0.621000 ;
        RECT 0.058000 0.399000 0.120000 0.494000 ;
        RECT 0.058000 0.399000 0.601000 0.454000 ;
        RECT 0.116000 0.386000 0.120000 0.494000 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.236000 0.539000 0.399000 0.627000 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.021000 0.550000 1.207000 0.645000 ;
        END
    END B0
    PIN C0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.769000 0.550000 0.905000 0.627000 ;
        RECT 1.282000 0.365000 1.407000 0.439000 ;
        RECT 1.345000 0.365000 1.407000 0.539000 ;
        RECT 0.843000 0.365000 0.905000 0.627000 ;
        RECT 0.843000 0.365000 1.407000 0.420000 ;
        END
    END C0
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 1.600000 1.280000 ;
        RECT 0.567000 0.925000 0.659000 1.280000 ;
        RECT 0.222000 0.925000 0.314000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 1.600000 0.080000 ;
        RECT 1.116000 -0.080000 1.208000 0.122000 ;
        RECT 0.407000 -0.080000 0.498000 0.122000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.323000 0.223000 1.414000 0.304000 ;
        RECT 1.086000 0.726000 1.177000 0.807000 ;
        RECT 0.762000 0.223000 0.980000 0.304000 ;
        RECT 0.051000 0.223000 0.143000 0.304000 ;
        RECT 1.100000 0.706000 1.177000 0.807000 ;
        RECT 0.749000 0.223000 0.980000 0.290000 ;
        RECT 1.471000 0.249000 1.533000 0.761000 ;
        RECT 1.323000 0.249000 1.533000 0.304000 ;
        RECT 1.100000 0.706000 1.533000 0.761000 ;
        RECT 0.051000 0.236000 1.414000 0.290000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 1.430000 0.881000 1.522000 0.962000 ;
        RECT 0.875000 0.688000 0.937000 0.949000 ;
        RECT 0.875000 0.894000 1.522000 0.949000 ;
        RECT 0.050000 0.688000 0.937000 0.743000 ;
    END
END AOI211X2

MACRO AND3X4
    CLASS CORE ;
    FOREIGN AND3X4 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 1.100000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.039000 0.433000 0.158000 0.577000 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.222000 0.560000 0.412000 0.633000 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.406000 0.433000 0.574000 0.500000 ;
        RECT 0.510000 0.433000 0.574000 0.576000 ;
        END
    END C
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 1.100000 1.280000 ;
        RECT 0.956000 0.933000 1.050000 1.280000 ;
        RECT 0.589000 0.908000 0.683000 1.280000 ;
        RECT 0.228000 0.908000 0.322000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 1.100000 0.080000 ;
        RECT 0.569000 -0.080000 0.664000 0.230000 ;
        RECT 0.956000 -0.080000 1.050000 0.122000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.956000 0.433000 1.061000 0.767000 ;
        RECT 0.956000 0.402000 1.040000 0.767000 ;
        RECT 0.792000 0.667000 1.061000 0.751000 ;
        RECT 0.765000 0.327000 0.829000 0.457000 ;
        RECT 0.765000 0.402000 1.040000 0.457000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 0.054000 0.257000 0.149000 0.338000 ;
        RECT 0.637000 0.317000 0.701000 0.802000 ;
        RECT 0.382000 0.270000 0.446000 0.371000 ;
        RECT 0.637000 0.546000 0.851000 0.601000 ;
        RECT 0.149000 0.270000 0.382000 0.325000 ;
        RECT 0.382000 0.317000 0.701000 0.371000 ;
        RECT 0.050000 0.748000 0.701000 0.802000 ;
    END
END AND3X4

MACRO AND3X2
    CLASS CORE ;
    FOREIGN AND3X2 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 0.900000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.038000 0.587000 0.142000 0.773000 ;
        RECT 0.038000 0.587000 0.155000 0.668000 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.218000 0.567000 0.342000 0.689000 ;
        RECT 0.280000 0.564000 0.342000 0.689000 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.447000 0.600000 0.540000 0.689000 ;
        RECT 0.398000 0.433000 0.510000 0.500000 ;
        RECT 0.447000 0.433000 0.510000 0.689000 ;
        END
    END C
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 0.900000 1.280000 ;
        RECT 0.545000 1.065000 0.638000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 0.900000 0.080000 ;
        RECT 0.507000 -0.080000 0.600000 0.122000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.715000 0.188000 0.807000 0.383000 ;
        RECT 0.753000 0.652000 0.845000 0.733000 ;
        RECT 0.768000 0.652000 0.845000 0.761000 ;
        RECT 0.715000 0.317000 0.845000 0.383000 ;
        RECT 0.783000 0.317000 0.845000 0.761000 ;
        RECT 0.783000 0.188000 0.807000 0.761000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 0.612000 0.488000 0.720000 0.583000 ;
        RECT 0.048000 0.954000 0.142000 1.049000 ;
        RECT 0.049000 0.298000 0.142000 0.379000 ;
        RECT 0.612000 0.488000 0.675000 0.829000 ;
        RECT 0.589000 0.324000 0.652000 0.543000 ;
        RECT 0.243000 0.774000 0.305000 1.008000 ;
        RECT 0.589000 0.488000 0.720000 0.543000 ;
        RECT 0.243000 0.774000 0.675000 0.829000 ;
        RECT 0.049000 0.324000 0.652000 0.379000 ;
        RECT 0.048000 0.954000 0.305000 1.008000 ;
        RECT 0.612000 0.324000 0.652000 0.829000 ;
    END
END AND3X2

MACRO AND2X4
    CLASS CORE ;
    FOREIGN AND2X4 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 0.900000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.038000 0.482000 0.142000 0.660000 ;
        RECT 0.038000 0.482000 0.145000 0.574000 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.218000 0.627000 0.322000 0.786000 ;
        RECT 0.312000 0.471000 0.375000 0.562000 ;
        RECT 0.259000 0.507000 0.322000 0.786000 ;
        RECT 0.259000 0.507000 0.375000 0.562000 ;
        RECT 0.312000 0.471000 0.322000 0.786000 ;
        END
    END B
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 0.900000 1.280000 ;
        RECT 0.046000 1.078000 0.146000 1.280000 ;
        RECT 0.755000 0.914000 0.848000 1.280000 ;
        RECT 0.394000 1.078000 0.487000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 0.900000 0.080000 ;
        RECT 0.755000 -0.080000 0.848000 0.243000 ;
        RECT 0.387000 -0.080000 0.480000 0.122000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.592000 0.326000 0.784000 0.433000 ;
        RECT 0.758000 0.433000 0.862000 0.767000 ;
        RECT 0.758000 0.331000 0.860000 0.798000 ;
        RECT 0.592000 0.331000 0.860000 0.433000 ;
        RECT 0.580000 0.717000 0.860000 0.798000 ;
        RECT 0.580000 0.717000 0.862000 0.767000 ;
        RECT 0.758000 0.326000 0.784000 0.798000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 0.440000 0.498000 0.663000 0.579000 ;
        RECT 0.049000 0.343000 0.142000 0.424000 ;
        RECT 0.440000 0.354000 0.503000 0.671000 ;
        RECT 0.386000 0.617000 0.449000 0.910000 ;
        RECT 0.202000 0.855000 0.449000 0.910000 ;
        RECT 0.386000 0.617000 0.503000 0.671000 ;
        RECT 0.202000 0.354000 0.503000 0.408000 ;
        RECT 0.142000 0.354000 0.440000 0.408000 ;
        RECT 0.049000 0.354000 0.386000 0.408000 ;
        RECT 0.440000 0.354000 0.449000 0.910000 ;
    END
END AND2X4

MACRO AND2X2
    CLASS CORE ;
    FOREIGN AND2X2 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 0.700000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.037000 0.504000 0.138000 0.633000 ;
        RECT 0.037000 0.504000 0.202000 0.585000 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.212000 0.833000 0.361000 0.935000 ;
        END
    END B
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 0.700000 1.280000 ;
        RECT 0.048000 1.078000 0.151000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 0.700000 0.080000 ;
        RECT 0.350000 -0.080000 0.440000 0.122000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.552000 0.227000 0.654000 0.390000 ;
        RECT 0.552000 0.688000 0.642000 1.002000 ;
        RECT 0.552000 0.195000 0.642000 0.390000 ;
        RECT 0.552000 0.688000 0.654000 0.767000 ;
        RECT 0.582000 0.227000 0.654000 0.439000 ;
        RECT 0.593000 0.227000 0.654000 0.767000 ;
        RECT 0.582000 0.195000 0.642000 0.439000 ;
        RECT 0.593000 0.195000 0.642000 1.002000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 0.216000 0.654000 0.325000 0.737000 ;
        RECT 0.264000 0.512000 0.521000 0.594000 ;
        RECT 0.048000 0.321000 0.138000 0.402000 ;
        RECT 0.264000 0.348000 0.325000 0.737000 ;
        RECT 0.048000 0.348000 0.325000 0.402000 ;
    END
END AND2X2

MACRO ADDHX2
    CLASS CORE ;
    FOREIGN ADDHX2 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 3.200000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 2.054000 0.454000 2.525000 0.535000 ;
        RECT 2.191000 0.439000 2.253000 0.535000 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.386000 0.438000 1.477000 0.519000 ;
        RECT 1.013000 0.538000 1.104000 0.619000 ;
        RECT 1.364000 0.438000 1.477000 0.506000 ;
        RECT 1.302000 0.439000 1.477000 0.506000 ;
        RECT 1.042000 0.451000 1.104000 0.619000 ;
        RECT 1.042000 0.451000 1.477000 0.506000 ;
        END
    END B
    PIN CO
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 2.890000 0.626000 2.982000 0.733000 ;
        RECT 2.902000 0.350000 2.985000 0.439000 ;
        RECT 2.964000 0.324000 3.099000 0.405000 ;
        RECT 2.902000 0.626000 2.967000 0.761000 ;
        RECT 2.902000 0.350000 2.964000 0.761000 ;
        RECT 2.902000 0.350000 3.099000 0.405000 ;
        RECT 2.964000 0.324000 2.985000 0.439000 ;
        END
    END CO
    PIN S
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.142000 0.674000 1.578000 0.755000 ;
        RECT 0.803000 0.306000 0.894000 0.387000 ;
        RECT 0.812000 0.687000 1.009000 0.761000 ;
        RECT 0.812000 0.687000 1.578000 0.755000 ;
        RECT 0.803000 0.306000 0.947000 0.374000 ;
        RECT 0.812000 0.669000 0.879000 0.761000 ;
        RECT 1.539000 0.306000 1.601000 0.392000 ;
        RECT 0.818000 0.306000 0.879000 0.761000 ;
        RECT 0.803000 0.319000 1.601000 0.374000 ;
        END
    END S
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 3.200000 1.280000 ;
        RECT 2.012000 1.002000 2.104000 1.280000 ;
        RECT 1.675000 1.065000 1.767000 1.280000 ;
        RECT 0.404000 1.078000 0.496000 1.280000 ;
        RECT 0.048000 1.002000 0.140000 1.280000 ;
        RECT 2.718000 0.989000 2.809000 1.280000 ;
        RECT 2.357000 0.989000 2.448000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 3.200000 0.080000 ;
        RECT 2.813000 -0.080000 2.905000 0.211000 ;
        RECT 2.474000 -0.080000 2.566000 0.220000 ;
        RECT 2.129000 -0.080000 2.221000 0.220000 ;
        RECT 0.404000 -0.080000 0.496000 0.122000 ;
        RECT 0.048000 -0.080000 0.140000 0.215000 ;
        END
    END VSS
    OBS
        LAYER Metal1 ;
        RECT 1.826000 0.604000 1.918000 0.762000 ;
        RECT 2.698000 0.514000 2.789000 0.595000 ;
        RECT 2.646000 0.313000 2.738000 0.394000 ;
        RECT 2.185000 0.713000 2.621000 0.794000 ;
        RECT 1.314000 0.969000 1.406000 1.050000 ;
        RECT 0.609000 0.652000 0.737000 0.733000 ;
        RECT 0.221000 0.652000 0.388000 0.733000 ;
        RECT 0.221000 0.325000 0.388000 0.406000 ;
        RECT 0.156000 0.505000 0.248000 0.586000 ;
        RECT 2.698000 0.514000 2.760000 0.658000 ;
        RECT 1.934000 0.158000 1.996000 0.379000 ;
        RECT 1.789000 0.289000 1.851000 0.658000 ;
        RECT 1.663000 0.158000 1.725000 0.896000 ;
        RECT 1.476000 0.842000 1.538000 1.024000 ;
        RECT 0.731000 0.843000 0.793000 0.939000 ;
        RECT 0.675000 0.302000 0.737000 0.733000 ;
        RECT 0.575000 0.952000 0.637000 1.050000 ;
        RECT 0.558000 0.158000 0.620000 0.248000 ;
        RECT 0.326000 0.193000 0.388000 0.898000 ;
        RECT 0.202000 0.850000 0.264000 1.007000 ;
        RECT 0.071000 0.531000 0.133000 0.905000 ;
        RECT 2.185000 0.713000 2.246000 0.896000 ;
        RECT 1.934000 0.324000 2.738000 0.379000 ;
        RECT 1.352000 0.158000 1.996000 0.213000 ;
        RECT 1.314000 0.969000 1.538000 1.024000 ;
        RECT 0.609000 0.302000 0.737000 0.357000 ;
        RECT 0.575000 0.995000 1.406000 1.050000 ;
        RECT 0.558000 0.158000 1.067000 0.213000 ;
        RECT 0.326000 0.843000 0.793000 0.898000 ;
        RECT 0.326000 0.193000 0.620000 0.248000 ;
        RECT 0.202000 0.952000 0.637000 1.007000 ;
        RECT 0.071000 0.850000 0.264000 0.905000 ;
        RECT 0.071000 0.531000 0.248000 0.586000 ;
        RECT 1.789000 0.604000 2.760000 0.658000 ;
        RECT 1.476000 0.842000 2.246000 0.896000 ;
        RECT 0.731000 0.885000 1.061000 0.939000 ;
        RECT 1.826000 0.289000 1.851000 0.762000 ;
    END
END ADDHX2

MACRO ADDFX2
    CLASS CORE ;
    FOREIGN ADDFX2 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 3.700000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.040000 0.560000 1.291000 0.640000 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.112000 0.486000 0.203000 0.567000 ;
        RECT 0.057000 0.512000 0.119000 0.627000 ;
        RECT 0.057000 0.512000 0.203000 0.567000 ;
        RECT 0.112000 0.486000 0.119000 0.627000 ;
        END
    END B
    PIN CI
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 2.296000 0.682000 2.461000 0.767000 ;
        RECT 2.400000 0.433000 2.461000 0.767000 ;
        RECT 2.400000 0.433000 2.532000 0.488000 ;
        END
    END CI
    PIN CO
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 3.078000 0.665000 3.199000 0.746000 ;
        RECT 3.078000 0.340000 3.205000 0.421000 ;
        RECT 3.078000 0.340000 3.139000 0.746000 ;
        RECT 3.053000 0.573000 3.139000 0.627000 ;
        END
    END CO
    PIN S
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 3.478000 0.306000 3.569000 0.424000 ;
        RECT 3.474000 0.665000 3.565000 0.746000 ;
        RECT 3.496000 0.306000 3.557000 0.746000 ;
        RECT 3.405000 0.306000 3.569000 0.361000 ;
        END
    END S
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 3.700000 1.280000 ;
        RECT 3.293000 1.078000 3.384000 1.280000 ;
        RECT 2.294000 1.078000 2.385000 1.280000 ;
        RECT 0.230000 1.078000 0.320000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 3.700000 0.080000 ;
        RECT 3.297000 -0.080000 3.388000 0.122000 ;
        RECT 2.600000 -0.080000 2.691000 0.122000 ;
        RECT 0.252000 -0.080000 0.343000 0.122000 ;
        RECT 1.171000 -0.080000 1.261000 0.199000 ;
        END
    END VSS
    OBS
        LAYER Metal1 ;
        RECT 1.479000 0.270000 1.570000 0.417000 ;
        RECT 0.048000 0.194000 0.139000 0.387000 ;
        RECT 1.403000 0.965000 1.785000 1.050000 ;
        RECT 1.353000 0.493000 1.658000 0.576000 ;
        RECT 2.892000 0.743000 2.983000 0.824000 ;
        RECT 2.700000 0.765000 2.791000 0.846000 ;
        RECT 2.226000 0.523000 2.339000 0.604000 ;
        RECT 1.719000 0.562000 1.850000 0.643000 ;
        RECT 1.531000 0.748000 1.622000 0.829000 ;
        RECT 0.402000 0.700000 0.531000 0.781000 ;
        RECT 0.307000 0.486000 0.398000 0.567000 ;
        RECT 0.048000 0.688000 0.330000 0.769000 ;
        RECT 1.723000 0.835000 1.814000 0.915000 ;
        RECT 1.478000 0.761000 1.622000 0.829000 ;
        RECT 0.268000 0.499000 0.398000 0.567000 ;
        RECT 1.531000 0.748000 1.648000 0.815000 ;
        RECT 2.728000 0.507000 2.790000 0.846000 ;
        RECT 2.473000 0.150000 2.535000 0.248000 ;
        RECT 2.226000 0.377000 2.288000 0.604000 ;
        RECT 2.158000 0.549000 2.220000 0.898000 ;
        RECT 2.034000 0.377000 2.096000 0.907000 ;
        RECT 1.911000 0.426000 1.973000 0.798000 ;
        RECT 1.723000 0.835000 1.785000 1.050000 ;
        RECT 1.719000 0.260000 1.781000 0.688000 ;
        RECT 1.508000 0.150000 1.570000 0.417000 ;
        RECT 1.353000 0.389000 1.415000 0.801000 ;
        RECT 0.734000 0.832000 0.796000 0.940000 ;
        RECT 0.715000 0.338000 0.777000 0.549000 ;
        RECT 0.268000 0.499000 0.330000 0.925000 ;
        RECT 3.373000 0.480000 3.434000 0.569000 ;
        RECT 3.280000 0.514000 3.341000 0.939000 ;
        RECT 2.910000 0.150000 2.971000 0.824000 ;
        RECT 2.787000 0.320000 2.848000 0.562000 ;
        RECT 2.730000 0.765000 2.791000 0.939000 ;
        RECT 2.595000 0.302000 2.656000 0.685000 ;
        RECT 2.523000 0.630000 2.584000 0.846000 ;
        RECT 2.447000 0.954000 2.508000 1.050000 ;
        RECT 2.351000 0.260000 2.412000 0.357000 ;
        RECT 2.036000 0.852000 2.097000 1.008000 ;
        RECT 1.842000 0.377000 1.903000 0.481000 ;
        RECT 1.753000 0.743000 1.814000 0.915000 ;
        RECT 1.587000 0.632000 1.648000 0.815000 ;
        RECT 1.478000 0.761000 1.539000 0.911000 ;
        RECT 1.048000 0.208000 1.109000 0.325000 ;
        RECT 0.980000 0.710000 1.041000 0.801000 ;
        RECT 0.925000 0.343000 0.986000 0.444000 ;
        RECT 0.857000 0.721000 0.918000 0.911000 ;
        RECT 0.788000 0.494000 0.849000 0.776000 ;
        RECT 0.638000 0.604000 0.699000 0.752000 ;
        RECT 0.593000 0.208000 0.654000 0.658000 ;
        RECT 0.506000 0.726000 0.567000 0.887000 ;
        RECT 0.470000 0.332000 0.531000 0.781000 ;
        RECT 0.382000 0.870000 0.443000 1.050000 ;
        RECT 0.307000 0.332000 0.368000 0.567000 ;
        RECT 2.730000 0.507000 2.790000 0.939000 ;
        RECT 2.036000 0.377000 2.096000 1.008000 ;
        RECT 1.587000 0.632000 1.781000 0.688000 ;
        RECT 3.280000 0.514000 3.434000 0.569000 ;
        RECT 2.910000 0.150000 3.013000 0.205000 ;
        RECT 2.728000 0.507000 2.848000 0.562000 ;
        RECT 2.523000 0.630000 2.656000 0.685000 ;
        RECT 2.473000 0.193000 2.971000 0.248000 ;
        RECT 2.447000 0.995000 3.034000 1.050000 ;
        RECT 2.351000 0.302000 2.656000 0.357000 ;
        RECT 2.158000 0.549000 2.339000 0.604000 ;
        RECT 1.915000 0.852000 2.097000 0.907000 ;
        RECT 1.842000 0.426000 1.973000 0.481000 ;
        RECT 1.753000 0.743000 1.973000 0.798000 ;
        RECT 1.508000 0.150000 2.535000 0.205000 ;
        RECT 1.048000 0.270000 1.570000 0.325000 ;
        RECT 0.980000 0.746000 1.415000 0.801000 ;
        RECT 0.925000 0.389000 1.415000 0.444000 ;
        RECT 0.857000 0.856000 1.539000 0.911000 ;
        RECT 0.788000 0.721000 0.918000 0.776000 ;
        RECT 0.715000 0.494000 0.849000 0.549000 ;
        RECT 0.593000 0.208000 1.109000 0.263000 ;
        RECT 0.506000 0.832000 0.796000 0.887000 ;
        RECT 0.402000 0.726000 0.567000 0.781000 ;
        RECT 0.382000 0.995000 1.785000 1.050000 ;
        RECT 0.268000 0.870000 0.443000 0.925000 ;
        RECT 0.048000 0.332000 0.368000 0.387000 ;
        RECT 2.730000 0.885000 3.341000 0.939000 ;
        RECT 2.036000 0.954000 2.508000 1.008000 ;
        RECT 1.719000 0.260000 2.412000 0.314000 ;
        RECT 1.478000 0.761000 1.648000 0.815000 ;
        RECT 0.593000 0.604000 0.699000 0.658000 ;
        RECT 1.587000 0.632000 1.622000 0.829000 ;
        RECT 1.753000 0.743000 1.785000 1.050000 ;
        RECT 0.506000 0.332000 0.531000 0.887000 ;
        RECT 0.307000 0.332000 0.330000 0.925000 ;
        RECT 0.638000 0.208000 0.654000 0.752000 ;
        RECT 1.531000 0.748000 1.539000 0.911000 ;
        RECT 2.787000 0.320000 2.790000 0.939000 ;
    END
END ADDFX2

MACRO ADDFHX2
    CLASS CORE ;
    FOREIGN ADDFHX2 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 5.900000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.191000 0.433000 0.327000 0.571000 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 3.363000 0.635000 3.699000 0.715000 ;
        RECT 3.527000 0.635000 3.588000 0.761000 ;
        END
    END B
    PIN CI
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 4.994000 0.546000 5.169000 0.649000 ;
        END
    END CI
    PIN CO
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 5.424000 0.331000 5.514000 0.412000 ;
        RECT 5.406000 0.344000 5.514000 0.412000 ;
        RECT 5.406000 0.344000 5.466000 0.761000 ;
        RECT 5.262000 0.706000 5.466000 0.761000 ;
        RECT 5.424000 0.331000 5.466000 0.761000 ;
        END
    END CO
    PIN S
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 5.737000 0.357000 5.845000 0.494000 ;
        RECT 5.755000 0.219000 5.845000 0.494000 ;
        RECT 5.723000 0.654000 5.812000 0.958000 ;
        RECT 5.737000 0.627000 5.812000 0.958000 ;
        RECT 5.737000 0.357000 5.797000 0.958000 ;
        RECT 5.755000 0.219000 5.797000 0.958000 ;
        END
    END S
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 5.900000 1.280000 ;
        RECT 4.834000 1.078000 4.940000 1.280000 ;
        RECT 5.533000 0.988000 5.623000 1.280000 ;
        RECT 3.615000 0.970000 3.705000 1.280000 ;
        RECT 5.202000 0.988000 5.291000 1.280000 ;
        RECT 3.237000 0.970000 3.326000 1.280000 ;
        RECT 0.873000 0.911000 0.962000 1.280000 ;
        RECT 0.291000 0.967000 0.380000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 5.900000 0.080000 ;
        RECT 5.224000 -0.080000 5.314000 0.122000 ;
        RECT 0.791000 -0.080000 0.881000 0.122000 ;
        RECT 0.260000 -0.080000 0.350000 0.122000 ;
        RECT 5.566000 -0.080000 5.655000 0.211000 ;
        RECT 3.481000 -0.080000 3.570000 0.122000 ;
        END
    END VSS
    OBS
        LAYER Metal1 ;
        RECT 0.047000 0.674000 0.137000 1.012000 ;
        RECT 4.450000 0.785000 4.539000 0.977000 ;
        RECT 4.261000 0.751000 4.350000 0.944000 ;
        RECT 4.028000 0.780000 4.117000 0.975000 ;
        RECT 3.805000 0.819000 3.894000 1.014000 ;
        RECT 3.426000 0.824000 3.515000 1.025000 ;
        RECT 4.776000 0.549000 4.888000 0.636000 ;
        RECT 1.387000 0.369000 1.470000 0.457000 ;
        RECT 4.639000 0.721000 4.729000 0.802000 ;
        RECT 3.681000 0.321000 3.770000 0.402000 ;
        RECT 1.625000 0.724000 1.714000 0.805000 ;
        RECT 1.441000 0.725000 1.530000 0.806000 ;
        RECT 0.770000 0.498000 0.860000 0.579000 ;
        RECT 0.644000 0.302000 0.734000 0.383000 ;
        RECT 0.460000 0.348000 0.550000 0.429000 ;
        RECT 0.394000 0.652000 0.484000 0.733000 ;
        RECT 0.047000 0.288000 0.137000 0.369000 ;
        RECT 4.042000 0.743000 4.117000 0.975000 ;
        RECT 2.546000 0.968000 2.621000 1.050000 ;
        RECT 1.058000 0.785000 1.156000 0.852000 ;
        RECT 0.678000 0.785000 0.776000 0.852000 ;
        RECT 3.983000 0.151000 4.048000 0.246000 ;
        RECT 5.278000 0.239000 5.339000 0.579000 ;
        RECT 4.827000 0.260000 4.888000 0.799000 ;
        RECT 4.464000 0.369000 4.525000 0.977000 ;
        RECT 4.275000 0.260000 4.336000 0.944000 ;
        RECT 3.987000 0.151000 4.048000 0.686000 ;
        RECT 3.866000 0.335000 3.927000 0.726000 ;
        RECT 3.745000 0.457000 3.806000 0.545000 ;
        RECT 3.290000 0.157000 3.351000 0.246000 ;
        RECT 2.901000 0.490000 2.962000 0.910000 ;
        RECT 2.721000 0.601000 2.782000 0.793000 ;
        RECT 2.612000 0.269000 2.673000 0.545000 ;
        RECT 2.491000 0.150000 2.552000 0.656000 ;
        RECT 1.739000 0.269000 1.800000 0.501000 ;
        RECT 1.409000 0.260000 1.470000 0.793000 ;
        RECT 1.095000 0.785000 1.156000 1.050000 ;
        RECT 0.933000 0.315000 0.994000 0.839000 ;
        RECT 0.456000 0.821000 0.517000 1.020000 ;
        RECT 0.423000 0.511000 0.484000 0.733000 ;
        RECT 0.076000 0.193000 0.137000 0.369000 ;
        RECT 5.527000 0.526000 5.587000 0.913000 ;
        RECT 4.950000 0.150000 5.010000 0.294000 ;
        RECT 4.654000 0.369000 4.714000 0.802000 ;
        RECT 4.123000 0.150000 4.183000 0.798000 ;
        RECT 3.819000 0.671000 3.879000 1.014000 ;
        RECT 3.426000 0.301000 3.486000 0.512000 ;
        RECT 3.146000 0.411000 3.206000 0.900000 ;
        RECT 3.146000 0.269000 3.206000 0.356000 ;
        RECT 3.025000 0.380000 3.085000 1.023000 ;
        RECT 2.356000 0.300000 2.416000 0.792000 ;
        RECT 2.118000 0.150000 2.178000 0.682000 ;
        RECT 1.951000 0.293000 2.011000 0.792000 ;
        RECT 1.929000 0.150000 1.989000 0.348000 ;
        RECT 1.829000 0.446000 1.889000 0.919000 ;
        RECT 1.625000 0.571000 1.685000 0.805000 ;
        RECT 1.549000 0.150000 1.609000 0.626000 ;
        RECT 1.266000 0.596000 1.326000 0.919000 ;
        RECT 1.195000 0.369000 1.255000 0.651000 ;
        RECT 1.065000 0.260000 1.125000 0.370000 ;
        RECT 0.943000 0.150000 1.003000 0.248000 ;
        RECT 0.475000 0.348000 0.535000 0.565000 ;
        RECT 0.062000 0.288000 0.122000 1.012000 ;
        RECT 4.950000 0.239000 5.339000 0.294000 ;
        RECT 4.827000 0.744000 5.092000 0.799000 ;
        RECT 4.827000 0.356000 5.114000 0.411000 ;
        RECT 4.654000 0.369000 4.767000 0.424000 ;
        RECT 4.464000 0.369000 4.576000 0.424000 ;
        RECT 4.450000 0.858000 5.587000 0.913000 ;
        RECT 4.123000 0.150000 5.010000 0.205000 ;
        RECT 4.042000 0.743000 4.183000 0.798000 ;
        RECT 3.426000 0.457000 3.806000 0.512000 ;
        RECT 3.146000 0.824000 3.894000 0.879000 ;
        RECT 3.146000 0.301000 3.486000 0.356000 ;
        RECT 2.733000 0.380000 3.085000 0.435000 ;
        RECT 2.721000 0.738000 2.836000 0.793000 ;
        RECT 2.612000 0.490000 2.962000 0.545000 ;
        RECT 2.612000 0.269000 3.206000 0.324000 ;
        RECT 2.546000 0.968000 3.085000 1.023000 ;
        RECT 2.491000 0.601000 2.782000 0.656000 ;
        RECT 2.491000 0.157000 3.351000 0.212000 ;
        RECT 2.293000 0.300000 2.416000 0.355000 ;
        RECT 2.118000 0.627000 2.293000 0.682000 ;
        RECT 2.118000 0.150000 2.552000 0.205000 ;
        RECT 1.951000 0.737000 2.493000 0.792000 ;
        RECT 1.829000 0.855000 2.962000 0.910000 ;
        RECT 1.739000 0.446000 1.889000 0.501000 ;
        RECT 1.549000 0.571000 1.685000 0.626000 ;
        RECT 1.266000 0.864000 1.889000 0.919000 ;
        RECT 1.195000 0.596000 1.326000 0.651000 ;
        RECT 1.095000 0.995000 2.621000 1.050000 ;
        RECT 0.943000 0.150000 1.989000 0.205000 ;
        RECT 0.644000 0.315000 1.125000 0.370000 ;
        RECT 0.456000 0.965000 0.631000 1.020000 ;
        RECT 0.076000 0.193000 1.003000 0.248000 ;
        RECT 0.047000 0.821000 0.517000 0.876000 ;
        RECT 4.275000 0.260000 4.888000 0.314000 ;
        RECT 3.681000 0.335000 3.927000 0.389000 ;
        RECT 3.290000 0.192000 4.048000 0.246000 ;
        RECT 3.146000 0.411000 3.360000 0.465000 ;
        RECT 1.065000 0.260000 1.470000 0.314000 ;
        RECT 0.678000 0.785000 1.156000 0.839000 ;
        RECT 0.423000 0.511000 0.860000 0.565000 ;
        RECT 0.076000 0.193000 0.122000 1.012000 ;
        RECT 1.951000 0.150000 1.989000 0.792000 ;
        RECT 1.441000 0.260000 1.470000 0.806000 ;
        RECT 3.866000 0.335000 3.879000 1.014000 ;
        RECT 0.475000 0.348000 0.484000 0.733000 ;
    END
END ADDFHX2

MACRO MX3X2
    CLASS CORE ;
    FOREIGN MX3X2 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 4.000000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 2.437000 0.525000 2.572000 0.633000 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.570000 0.433000 1.702000 0.540000 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.037000 0.433000 0.200000 0.549000 ;
        RECT 0.111000 0.433000 0.200000 0.550000 ;
        END
    END C
    PIN S0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.524000 0.960000 0.614000 1.040000 ;
        RECT 0.524000 0.960000 0.639000 1.027000 ;
        RECT 0.626000 0.951000 0.752000 1.014000 ;
        RECT 2.012000 0.951000 2.072000 1.033000 ;
        RECT 0.626000 0.951000 2.072000 1.006000 ;
        RECT 0.524000 0.960000 0.752000 1.014000 ;
        RECT 0.626000 0.951000 0.639000 1.027000 ;
        END
    END S0
    PIN S1
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 3.348000 0.579000 3.491000 0.660000 ;
        RECT 2.819000 0.839000 2.920000 0.919000 ;
        RECT 3.348000 0.579000 3.408000 0.894000 ;
        RECT 2.819000 0.839000 3.408000 0.894000 ;
        END
    END S1
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 4.000000 1.280000 ;
        RECT 3.611000 0.877000 3.701000 1.280000 ;
        RECT 0.047000 0.757000 0.137000 1.280000 ;
        RECT 2.501000 1.078000 2.590000 1.280000 ;
        RECT 1.510000 1.078000 1.599000 1.280000 ;
        RECT 1.016000 1.078000 1.105000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 4.000000 0.080000 ;
        RECT 3.611000 -0.080000 3.701000 0.210000 ;
        RECT 2.502000 -0.080000 2.592000 0.122000 ;
        RECT 0.047000 -0.080000 0.137000 0.364000 ;
        RECT 1.510000 -0.080000 1.599000 0.122000 ;
        RECT 1.049000 -0.080000 1.138000 0.122000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 3.817000 0.701000 3.906000 1.006000 ;
        RECT 3.817000 0.180000 3.906000 0.373000 ;
        RECT 3.846000 0.180000 3.906000 1.006000 ;
        RECT 3.817000 0.706000 3.943000 0.761000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 2.080000 0.206000 2.190000 0.310000 ;
        RECT 2.088000 0.200000 2.190000 0.310000 ;
        RECT 2.997000 0.200000 3.087000 0.402000 ;
        RECT 2.295000 0.692000 2.385000 0.885000 ;
        RECT 0.751000 0.171000 0.841000 0.261000 ;
        RECT 0.428000 0.186000 0.518000 0.379000 ;
        RECT 0.237000 0.742000 0.327000 0.965000 ;
        RECT 0.237000 0.186000 0.327000 0.379000 ;
        RECT 3.427000 0.157000 3.516000 0.350000 ;
        RECT 3.207000 0.194000 3.296000 0.492000 ;
        RECT 3.507000 0.408000 3.593000 0.508000 ;
        RECT 3.115000 0.681000 3.204000 0.762000 ;
        RECT 2.925000 0.681000 3.014000 0.762000 ;
        RECT 2.702000 0.688000 2.792000 0.769000 ;
        RECT 2.702000 0.336000 2.931000 0.417000 ;
        RECT 2.295000 0.317000 2.385000 0.398000 ;
        RECT 2.066000 0.679000 2.155000 0.760000 ;
        RECT 1.808000 0.329000 2.004000 0.410000 ;
        RECT 1.792000 0.526000 1.881000 0.607000 ;
        RECT 1.710000 0.705000 1.800000 0.786000 ;
        RECT 1.231000 0.689000 1.320000 0.770000 ;
        RECT 0.812000 0.679000 0.901000 0.760000 ;
        RECT 0.730000 0.524000 0.866000 0.605000 ;
        RECT 0.606000 0.325000 0.743000 0.406000 ;
        RECT 0.427000 0.814000 0.516000 0.895000 ;
        RECT 1.260000 0.346000 1.340000 0.650000 ;
        RECT 1.792000 0.526000 1.867000 0.650000 ;
        RECT 1.244000 0.346000 1.340000 0.411000 ;
        RECT 2.997000 0.200000 3.058000 0.592000 ;
        RECT 2.939000 0.537000 3.000000 0.762000 ;
        RECT 2.295000 0.317000 2.356000 0.885000 ;
        RECT 2.080000 0.206000 2.141000 0.760000 ;
        RECT 1.943000 0.329000 2.004000 0.773000 ;
        RECT 1.751000 0.150000 1.812000 0.261000 ;
        RECT 0.805000 0.346000 0.866000 0.605000 ;
        RECT 0.606000 0.325000 0.667000 0.746000 ;
        RECT 0.266000 0.186000 0.327000 0.965000 ;
        RECT 3.659000 0.295000 3.719000 0.787000 ;
        RECT 3.472000 0.732000 3.532000 1.042000 ;
        RECT 3.144000 0.437000 3.204000 0.762000 ;
        RECT 2.717000 0.336000 2.777000 0.769000 ;
        RECT 2.667000 0.939000 2.727000 1.042000 ;
        RECT 2.157000 0.842000 2.217000 0.994000 ;
        RECT 1.497000 0.825000 1.557000 0.896000 ;
        RECT 1.260000 0.346000 1.320000 0.770000 ;
        RECT 1.107000 0.814000 1.167000 0.880000 ;
        RECT 0.447000 0.186000 0.507000 0.895000 ;
        RECT 3.472000 0.732000 3.719000 0.787000 ;
        RECT 3.427000 0.295000 3.719000 0.350000 ;
        RECT 3.144000 0.437000 3.593000 0.492000 ;
        RECT 2.939000 0.537000 3.058000 0.592000 ;
        RECT 2.667000 0.987000 3.532000 1.042000 ;
        RECT 2.157000 0.939000 2.727000 0.994000 ;
        RECT 2.088000 0.200000 3.087000 0.255000 ;
        RECT 1.751000 0.150000 1.897000 0.205000 ;
        RECT 1.710000 0.718000 2.004000 0.773000 ;
        RECT 1.260000 0.595000 1.867000 0.650000 ;
        RECT 1.107000 0.825000 1.557000 0.880000 ;
        RECT 0.805000 0.346000 1.340000 0.401000 ;
        RECT 0.751000 0.206000 1.812000 0.261000 ;
        RECT 0.427000 0.814000 1.167000 0.869000 ;
        RECT 1.497000 0.842000 2.217000 0.896000 ;
        RECT 0.606000 0.692000 0.901000 0.746000 ;
        RECT 2.088000 0.200000 2.141000 0.760000 ;
        RECT 2.997000 0.200000 3.000000 0.762000 ;
    END
END MX3X2

MACRO TLATNTSCAX2
    CLASS CORE ;
    FOREIGN TLATNTSCAX2 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 3.300000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER Metal1 ;
        RECT 2.992000 0.433000 3.089000 0.580000 ;
        END
    END CK
    PIN E
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 2.816000 0.504000 2.916000 0.654000 ;
        END
    END E
    PIN ECK
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 2.342000 0.669000 2.432000 0.761000 ;
        RECT 2.342000 0.338000 2.432000 0.419000 ;
        RECT 2.342000 0.627000 2.412000 0.761000 ;
        RECT 2.351000 0.338000 2.412000 0.761000 ;
        RECT 2.314000 0.706000 2.432000 0.761000 ;
        END
    END ECK
    PIN SE
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.824000 0.464000 1.037000 0.545000 ;
        RECT 0.925000 0.439000 0.986000 0.545000 ;
        END
    END SE
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 3.300000 1.280000 ;
        RECT 0.884000 1.002000 0.976000 1.280000 ;
        RECT 1.963000 0.839000 2.053000 1.280000 ;
        RECT 1.384000 1.078000 1.474000 1.280000 ;
        RECT 0.247000 1.078000 0.337000 1.280000 ;
        RECT 2.937000 0.733000 3.026000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 3.300000 0.080000 ;
        RECT 0.884000 -0.080000 0.976000 0.200000 ;
        RECT 2.937000 -0.080000 3.026000 0.122000 ;
        RECT 1.953000 -0.080000 2.042000 0.122000 ;
        RECT 1.529000 -0.080000 1.618000 0.122000 ;
        RECT 0.258000 -0.080000 0.347000 0.122000 ;
        END
    END VSS
    OBS
        LAYER Metal1 ;
        RECT 1.126000 0.477000 1.226000 0.655000 ;
        RECT 0.405000 0.574000 0.500000 0.773000 ;
        RECT 0.546000 0.844000 0.638000 0.939000 ;
        RECT 1.126000 0.464000 1.216000 0.655000 ;
        RECT 0.032000 0.954000 0.137000 1.042000 ;
        RECT 0.304000 0.313000 0.480000 0.395000 ;
        RECT 3.126000 0.752000 3.216000 0.833000 ;
        RECT 3.095000 0.298000 3.184000 0.379000 ;
        RECT 2.737000 0.343000 2.826000 0.424000 ;
        RECT 2.686000 0.769000 2.826000 0.850000 ;
        RECT 2.671000 0.955000 2.761000 1.036000 ;
        RECT 2.532000 0.813000 2.621000 0.894000 ;
        RECT 2.532000 0.338000 2.621000 0.419000 ;
        RECT 2.153000 0.813000 2.242000 0.894000 ;
        RECT 2.153000 0.338000 2.242000 0.419000 ;
        RECT 1.880000 0.490000 2.093000 0.571000 ;
        RECT 1.753000 0.312000 1.842000 0.393000 ;
        RECT 1.539000 0.952000 1.629000 1.033000 ;
        RECT 1.384000 0.736000 1.474000 0.817000 ;
        RECT 1.332000 0.150000 1.421000 0.231000 ;
        RECT 1.224000 0.300000 1.313000 0.381000 ;
        RECT 1.661000 0.490000 2.093000 0.558000 ;
        RECT 1.332000 0.163000 1.447000 0.231000 ;
        RECT 3.095000 0.312000 3.213000 0.379000 ;
        RECT 1.537000 0.612000 1.600000 0.694000 ;
        RECT 1.537000 0.600000 1.599000 0.694000 ;
        RECT 2.546000 0.338000 2.607000 0.894000 ;
        RECT 2.153000 0.710000 2.214000 0.894000 ;
        RECT 1.788000 0.710000 1.849000 0.890000 ;
        RECT 1.550000 0.313000 1.611000 0.545000 ;
        RECT 1.539000 0.877000 1.600000 1.033000 ;
        RECT 1.050000 0.176000 1.111000 0.325000 ;
        RECT 0.759000 0.877000 0.820000 1.050000 ;
        RECT 0.417000 0.161000 0.478000 0.248000 ;
        RECT 3.153000 0.312000 3.213000 0.833000 ;
        RECT 3.095000 0.193000 3.155000 0.379000 ;
        RECT 2.686000 0.369000 2.746000 1.036000 ;
        RECT 2.154000 0.338000 2.214000 0.894000 ;
        RECT 1.661000 0.490000 1.721000 0.817000 ;
        RECT 1.387000 0.163000 1.447000 0.248000 ;
        RECT 0.662000 0.443000 0.722000 0.655000 ;
        RECT 0.595000 0.749000 0.655000 0.899000 ;
        RECT 0.541000 0.270000 0.601000 0.518000 ;
        RECT 0.404000 0.954000 0.464000 1.050000 ;
        RECT 0.304000 0.313000 0.364000 0.629000 ;
        RECT 0.183000 0.193000 0.243000 0.348000 ;
        RECT 0.153000 0.293000 0.213000 0.899000 ;
        RECT 0.062000 0.150000 0.122000 0.233000 ;
        RECT 0.032000 0.179000 0.092000 1.042000 ;
        RECT 2.686000 0.369000 2.826000 0.424000 ;
        RECT 2.153000 0.839000 2.621000 0.894000 ;
        RECT 1.753000 0.338000 2.242000 0.393000 ;
        RECT 1.550000 0.490000 2.093000 0.545000 ;
        RECT 1.387000 0.193000 3.155000 0.248000 ;
        RECT 1.384000 0.762000 1.721000 0.817000 ;
        RECT 1.332000 0.313000 1.611000 0.368000 ;
        RECT 1.313000 0.313000 1.550000 0.368000 ;
        RECT 1.224000 0.313000 1.539000 0.368000 ;
        RECT 1.050000 0.176000 1.447000 0.231000 ;
        RECT 0.759000 0.877000 1.600000 0.932000 ;
        RECT 0.662000 0.600000 1.599000 0.655000 ;
        RECT 0.595000 0.749000 1.474000 0.804000 ;
        RECT 0.541000 0.270000 1.111000 0.325000 ;
        RECT 0.425000 0.463000 0.601000 0.518000 ;
        RECT 0.404000 0.995000 0.820000 1.050000 ;
        RECT 0.304000 0.574000 0.722000 0.629000 ;
        RECT 0.183000 0.193000 0.478000 0.248000 ;
        RECT 0.153000 0.844000 0.655000 0.899000 ;
        RECT 0.153000 0.293000 0.243000 0.348000 ;
        RECT 1.788000 0.710000 2.214000 0.764000 ;
        RECT 0.417000 0.161000 0.638000 0.215000 ;
        RECT 0.122000 0.954000 0.464000 1.008000 ;
        RECT 0.032000 0.954000 0.364000 1.008000 ;
        RECT 0.032000 0.179000 0.122000 0.233000 ;
        RECT 0.595000 0.749000 0.638000 0.939000 ;
        RECT 1.387000 0.150000 1.421000 0.248000 ;
        RECT 0.183000 0.193000 0.213000 0.899000 ;
        RECT 0.062000 0.150000 0.092000 1.042000 ;
        RECT 3.155000 0.298000 3.184000 0.833000 ;
        RECT 2.737000 0.343000 2.746000 1.036000 ;
        RECT 3.153000 0.193000 3.155000 0.833000 ;
    END
END TLATNTSCAX2

MACRO BUFX6
    CLASS CORE ;
    FOREIGN BUFX6 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 1.300000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.160000 0.474000 0.391000 0.555000 ;
        RECT 0.246000 0.439000 0.311000 0.555000 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 1.300000 1.280000 ;
        RECT 0.422000 1.078000 0.518000 1.280000 ;
        RECT 1.154000 0.877000 1.249000 1.280000 ;
        RECT 0.794000 0.877000 0.889000 1.280000 ;
        RECT 0.051000 0.844000 0.146000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 1.300000 0.080000 ;
        RECT 0.816000 -0.080000 0.912000 0.215000 ;
        RECT 0.456000 -0.080000 0.552000 0.215000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.803000 0.433000 1.240000 0.767000 ;
        RECT 0.803000 0.321000 1.126000 0.767000 ;
        RECT 0.782000 0.625000 1.240000 0.757000 ;
        RECT 0.782000 0.321000 1.126000 0.440000 ;
        RECT 0.636000 0.321000 1.126000 0.402000 ;
        RECT 0.613000 0.676000 1.240000 0.757000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 0.484000 0.519000 0.718000 0.600000 ;
        RECT 0.253000 0.274000 0.349000 0.355000 ;
        RECT 0.231000 0.657000 0.326000 0.738000 ;
        RECT 0.484000 0.300000 0.549000 0.712000 ;
        RECT 0.253000 0.300000 0.549000 0.355000 ;
        RECT 0.231000 0.657000 0.549000 0.712000 ;
    END
END BUFX6

MACRO MEM1
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN MEM1 0 0 ;
  SIZE 426.965 BY 114.215 ;
  SYMMETRY X Y R90 ;
  PIN A[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12.00 77.64 12.66 78.30 ;
      LAYER Metal6 ;
        RECT 12.00 77.64 12.66 78.30 ;
      LAYER Metal3 ;
        RECT 12.00 77.64 12.66 78.30 ;
      LAYER Metal4 ;
        RECT 12.00 77.64 12.66 78.30 ;
    END
  END A[0]
  PIN A[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12.00 71.52 12.66 72.18 ;
      LAYER Metal6 ;
        RECT 12.00 71.52 12.66 72.18 ;
      LAYER Metal3 ;
        RECT 12.00 71.52 12.66 72.18 ;
      LAYER Metal4 ;
        RECT 12.00 71.52 12.66 72.18 ;
    END
  END A[1]
  PIN A[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12.00 68.42 12.66 69.08 ;
      LAYER Metal6 ;
        RECT 12.00 68.42 12.66 69.08 ;
      LAYER Metal3 ;
        RECT 12.00 68.42 12.66 69.08 ;
      LAYER Metal4 ;
        RECT 12.00 68.42 12.66 69.08 ;
    END
  END A[2]
  PIN A[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12.00 62.30 12.66 62.96 ;
      LAYER Metal6 ;
        RECT 12.00 62.30 12.66 62.96 ;
      LAYER Metal3 ;
        RECT 12.00 62.30 12.66 62.96 ;
      LAYER Metal4 ;
        RECT 12.00 62.30 12.66 62.96 ;
    END
  END A[3]
  PIN A[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12.00 59.28 12.66 59.94 ;
      LAYER Metal6 ;
        RECT 12.00 59.28 12.66 59.94 ;
      LAYER Metal3 ;
        RECT 12.00 59.28 12.66 59.94 ;
      LAYER Metal4 ;
        RECT 12.00 59.28 12.66 59.94 ;
    END
  END A[4]
  PIN A[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12.00 56.18 12.66 56.84 ;
      LAYER Metal6 ;
        RECT 12.00 56.18 12.66 56.84 ;
      LAYER Metal3 ;
        RECT 12.00 56.18 12.66 56.84 ;
      LAYER Metal4 ;
        RECT 12.00 56.18 12.66 56.84 ;
    END
  END A[5]
  PIN A[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12.00 50.06 12.66 50.72 ;
      LAYER Metal6 ;
        RECT 12.00 50.06 12.66 50.72 ;
      LAYER Metal3 ;
        RECT 12.00 50.06 12.66 50.72 ;
      LAYER Metal4 ;
        RECT 12.00 50.06 12.66 50.72 ;
    END
  END A[6]
  PIN A[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12.00 47.04 12.66 47.70 ;
      LAYER Metal6 ;
        RECT 12.00 47.04 12.66 47.70 ;
      LAYER Metal3 ;
        RECT 12.00 47.04 12.66 47.70 ;
      LAYER Metal4 ;
        RECT 12.00 47.04 12.66 47.70 ;
    END
  END A[7]
  PIN CE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 228.44 12.00 229.09 12.66 ;
      LAYER Metal6 ;
        RECT 228.44 12.00 229.09 12.66 ;
      LAYER Metal3 ;
        RECT 228.44 12.00 229.09 12.66 ;
      LAYER Metal4 ;
        RECT 228.44 12.00 229.09 12.66 ;
    END
  END CE
  PIN CK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER Metal5 ;
        RECT 238.18 12.00 238.84 12.66 ;
      LAYER Metal6 ;
        RECT 238.18 12.00 238.84 12.66 ;
      LAYER Metal3 ;
        RECT 238.18 12.00 238.84 12.66 ;
      LAYER Metal4 ;
        RECT 238.18 12.00 238.84 12.66 ;
    END
  END CK
  PIN D[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 20.48 12.00 21.14 12.66 ;
      LAYER Metal6 ;
        RECT 20.48 12.00 21.14 12.66 ;
      LAYER Metal3 ;
        RECT 20.48 12.00 21.14 12.66 ;
      LAYER Metal4 ;
        RECT 20.48 12.00 21.14 12.66 ;
    END
  END D[0]
  PIN D[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 129.00 12.00 129.66 12.66 ;
      LAYER Metal6 ;
        RECT 129.00 12.00 129.66 12.66 ;
      LAYER Metal3 ;
        RECT 129.00 12.00 129.66 12.66 ;
      LAYER Metal4 ;
        RECT 129.00 12.00 129.66 12.66 ;
    END
  END D[10]
  PIN D[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 137.04 12.00 137.70 12.66 ;
      LAYER Metal6 ;
        RECT 137.04 12.00 137.70 12.66 ;
      LAYER Metal3 ;
        RECT 137.04 12.00 137.70 12.66 ;
      LAYER Metal4 ;
        RECT 137.04 12.00 137.70 12.66 ;
    END
  END D[11]
  PIN D[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 151.34 12.00 152.00 12.66 ;
      LAYER Metal6 ;
        RECT 151.34 12.00 152.00 12.66 ;
      LAYER Metal3 ;
        RECT 151.34 12.00 152.00 12.66 ;
      LAYER Metal4 ;
        RECT 151.34 12.00 152.00 12.66 ;
    END
  END D[12]
  PIN D[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 159.38 12.00 160.04 12.66 ;
      LAYER Metal6 ;
        RECT 159.38 12.00 160.04 12.66 ;
      LAYER Metal3 ;
        RECT 159.38 12.00 160.04 12.66 ;
      LAYER Metal4 ;
        RECT 159.38 12.00 160.04 12.66 ;
    END
  END D[13]
  PIN D[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 172.62 12.00 173.28 12.66 ;
      LAYER Metal6 ;
        RECT 172.62 12.00 173.28 12.66 ;
      LAYER Metal3 ;
        RECT 172.62 12.00 173.28 12.66 ;
      LAYER Metal4 ;
        RECT 172.62 12.00 173.28 12.66 ;
    END
  END D[14]
  PIN D[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 180.66 12.00 181.32 12.66 ;
      LAYER Metal6 ;
        RECT 180.66 12.00 181.32 12.66 ;
      LAYER Metal3 ;
        RECT 180.66 12.00 181.32 12.66 ;
      LAYER Metal4 ;
        RECT 180.66 12.00 181.32 12.66 ;
    END
  END D[15]
  PIN D[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 245.65 12.00 246.31 12.66 ;
      LAYER Metal6 ;
        RECT 245.65 12.00 246.31 12.66 ;
      LAYER Metal3 ;
        RECT 245.65 12.00 246.31 12.66 ;
      LAYER Metal4 ;
        RECT 245.65 12.00 246.31 12.66 ;
    END
  END D[16]
  PIN D[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 253.69 12.00 254.34 12.66 ;
      LAYER Metal6 ;
        RECT 253.69 12.00 254.34 12.66 ;
      LAYER Metal3 ;
        RECT 253.69 12.00 254.34 12.66 ;
      LAYER Metal4 ;
        RECT 253.69 12.00 254.34 12.66 ;
    END
  END D[17]
  PIN D[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 266.93 12.00 267.58 12.66 ;
      LAYER Metal6 ;
        RECT 266.93 12.00 267.58 12.66 ;
      LAYER Metal3 ;
        RECT 266.93 12.00 267.58 12.66 ;
      LAYER Metal4 ;
        RECT 266.93 12.00 267.58 12.66 ;
    END
  END D[18]
  PIN D[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 274.96 12.00 275.62 12.66 ;
      LAYER Metal6 ;
        RECT 274.96 12.00 275.62 12.66 ;
      LAYER Metal3 ;
        RECT 274.96 12.00 275.62 12.66 ;
      LAYER Metal4 ;
        RECT 274.96 12.00 275.62 12.66 ;
    END
  END D[19]
  PIN D[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 28.52 12.00 29.18 12.66 ;
      LAYER Metal6 ;
        RECT 28.52 12.00 29.18 12.66 ;
      LAYER Metal3 ;
        RECT 28.52 12.00 29.18 12.66 ;
      LAYER Metal4 ;
        RECT 28.52 12.00 29.18 12.66 ;
    END
  END D[1]
  PIN D[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 289.26 12.00 289.93 12.66 ;
      LAYER Metal6 ;
        RECT 289.26 12.00 289.93 12.66 ;
      LAYER Metal3 ;
        RECT 289.26 12.00 289.93 12.66 ;
      LAYER Metal4 ;
        RECT 289.26 12.00 289.93 12.66 ;
    END
  END D[20]
  PIN D[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 297.31 12.00 297.96 12.66 ;
      LAYER Metal6 ;
        RECT 297.31 12.00 297.96 12.66 ;
      LAYER Metal3 ;
        RECT 297.31 12.00 297.96 12.66 ;
      LAYER Metal4 ;
        RECT 297.31 12.00 297.96 12.66 ;
    END
  END D[21]
  PIN D[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 310.55 12.00 311.20 12.66 ;
      LAYER Metal6 ;
        RECT 310.55 12.00 311.20 12.66 ;
      LAYER Metal3 ;
        RECT 310.55 12.00 311.20 12.66 ;
      LAYER Metal4 ;
        RECT 310.55 12.00 311.20 12.66 ;
    END
  END D[22]
  PIN D[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 318.58 12.00 319.25 12.66 ;
      LAYER Metal6 ;
        RECT 318.58 12.00 319.25 12.66 ;
      LAYER Metal3 ;
        RECT 318.58 12.00 319.25 12.66 ;
      LAYER Metal4 ;
        RECT 318.58 12.00 319.25 12.66 ;
    END
  END D[23]
  PIN D[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 332.88 12.00 333.55 12.66 ;
      LAYER Metal6 ;
        RECT 332.88 12.00 333.55 12.66 ;
      LAYER Metal3 ;
        RECT 332.88 12.00 333.55 12.66 ;
      LAYER Metal4 ;
        RECT 332.88 12.00 333.55 12.66 ;
    END
  END D[24]
  PIN D[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 340.93 12.00 341.58 12.66 ;
      LAYER Metal6 ;
        RECT 340.93 12.00 341.58 12.66 ;
      LAYER Metal3 ;
        RECT 340.93 12.00 341.58 12.66 ;
      LAYER Metal4 ;
        RECT 340.93 12.00 341.58 12.66 ;
    END
  END D[25]
  PIN D[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 354.17 12.00 354.82 12.66 ;
      LAYER Metal6 ;
        RECT 354.17 12.00 354.82 12.66 ;
      LAYER Metal3 ;
        RECT 354.17 12.00 354.82 12.66 ;
      LAYER Metal4 ;
        RECT 354.17 12.00 354.82 12.66 ;
    END
  END D[26]
  PIN D[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 362.20 12.00 362.87 12.66 ;
      LAYER Metal6 ;
        RECT 362.20 12.00 362.87 12.66 ;
      LAYER Metal3 ;
        RECT 362.20 12.00 362.87 12.66 ;
      LAYER Metal4 ;
        RECT 362.20 12.00 362.87 12.66 ;
    END
  END D[27]
  PIN D[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 376.50 12.00 377.17 12.66 ;
      LAYER Metal6 ;
        RECT 376.50 12.00 377.17 12.66 ;
      LAYER Metal3 ;
        RECT 376.50 12.00 377.17 12.66 ;
      LAYER Metal4 ;
        RECT 376.50 12.00 377.17 12.66 ;
    END
  END D[28]
  PIN D[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 384.55 12.00 385.20 12.66 ;
      LAYER Metal6 ;
        RECT 384.55 12.00 385.20 12.66 ;
      LAYER Metal3 ;
        RECT 384.55 12.00 385.20 12.66 ;
      LAYER Metal4 ;
        RECT 384.55 12.00 385.20 12.66 ;
    END
  END D[29]
  PIN D[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 41.76 12.00 42.42 12.66 ;
      LAYER Metal6 ;
        RECT 41.76 12.00 42.42 12.66 ;
      LAYER Metal3 ;
        RECT 41.76 12.00 42.42 12.66 ;
      LAYER Metal4 ;
        RECT 41.76 12.00 42.42 12.66 ;
    END
  END D[2]
  PIN D[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 397.79 12.00 398.44 12.66 ;
      LAYER Metal6 ;
        RECT 397.79 12.00 398.44 12.66 ;
      LAYER Metal3 ;
        RECT 397.79 12.00 398.44 12.66 ;
      LAYER Metal4 ;
        RECT 397.79 12.00 398.44 12.66 ;
    END
  END D[30]
  PIN D[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 405.82 12.00 406.49 12.66 ;
      LAYER Metal6 ;
        RECT 405.82 12.00 406.49 12.66 ;
      LAYER Metal3 ;
        RECT 405.82 12.00 406.49 12.66 ;
      LAYER Metal4 ;
        RECT 405.82 12.00 406.49 12.66 ;
    END
  END D[31]
  PIN D[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 49.80 12.00 50.46 12.66 ;
      LAYER Metal6 ;
        RECT 49.80 12.00 50.46 12.66 ;
      LAYER Metal3 ;
        RECT 49.80 12.00 50.46 12.66 ;
      LAYER Metal4 ;
        RECT 49.80 12.00 50.46 12.66 ;
    END
  END D[3]
  PIN D[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 64.10 12.00 64.76 12.66 ;
      LAYER Metal6 ;
        RECT 64.10 12.00 64.76 12.66 ;
      LAYER Metal3 ;
        RECT 64.10 12.00 64.76 12.66 ;
      LAYER Metal4 ;
        RECT 64.10 12.00 64.76 12.66 ;
    END
  END D[4]
  PIN D[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 72.14 12.00 72.80 12.66 ;
      LAYER Metal6 ;
        RECT 72.14 12.00 72.80 12.66 ;
      LAYER Metal3 ;
        RECT 72.14 12.00 72.80 12.66 ;
      LAYER Metal4 ;
        RECT 72.14 12.00 72.80 12.66 ;
    END
  END D[5]
  PIN D[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 85.38 12.00 86.04 12.66 ;
      LAYER Metal6 ;
        RECT 85.38 12.00 86.04 12.66 ;
      LAYER Metal3 ;
        RECT 85.38 12.00 86.04 12.66 ;
      LAYER Metal4 ;
        RECT 85.38 12.00 86.04 12.66 ;
    END
  END D[6]
  PIN D[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 93.42 12.00 94.08 12.66 ;
      LAYER Metal6 ;
        RECT 93.42 12.00 94.08 12.66 ;
      LAYER Metal3 ;
        RECT 93.42 12.00 94.08 12.66 ;
      LAYER Metal4 ;
        RECT 93.42 12.00 94.08 12.66 ;
    END
  END D[7]
  PIN D[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 107.72 12.00 108.38 12.66 ;
      LAYER Metal6 ;
        RECT 107.72 12.00 108.38 12.66 ;
      LAYER Metal3 ;
        RECT 107.72 12.00 108.38 12.66 ;
      LAYER Metal4 ;
        RECT 107.72 12.00 108.38 12.66 ;
    END
  END D[8]
  PIN D[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 115.76 12.00 116.42 12.66 ;
      LAYER Metal6 ;
        RECT 115.76 12.00 116.42 12.66 ;
      LAYER Metal3 ;
        RECT 115.76 12.00 116.42 12.66 ;
      LAYER Metal4 ;
        RECT 115.76 12.00 116.42 12.66 ;
    END
  END D[9]
  PIN Q[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 23.06 12.00 23.72 12.66 ;
      LAYER Metal6 ;
        RECT 23.06 12.00 23.72 12.66 ;
      LAYER Metal3 ;
        RECT 23.06 12.00 23.72 12.66 ;
      LAYER Metal4 ;
        RECT 23.06 12.00 23.72 12.66 ;
    END
  END Q[0]
  PIN Q[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 131.58 12.00 132.24 12.66 ;
      LAYER Metal6 ;
        RECT 131.58 12.00 132.24 12.66 ;
      LAYER Metal3 ;
        RECT 131.58 12.00 132.24 12.66 ;
      LAYER Metal4 ;
        RECT 131.58 12.00 132.24 12.66 ;
    END
  END Q[10]
  PIN Q[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 134.46 12.00 135.12 12.66 ;
      LAYER Metal6 ;
        RECT 134.46 12.00 135.12 12.66 ;
      LAYER Metal3 ;
        RECT 134.46 12.00 135.12 12.66 ;
      LAYER Metal4 ;
        RECT 134.46 12.00 135.12 12.66 ;
    END
  END Q[11]
  PIN Q[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 153.92 12.00 154.58 12.66 ;
      LAYER Metal6 ;
        RECT 153.92 12.00 154.58 12.66 ;
      LAYER Metal3 ;
        RECT 153.92 12.00 154.58 12.66 ;
      LAYER Metal4 ;
        RECT 153.92 12.00 154.58 12.66 ;
    END
  END Q[12]
  PIN Q[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 156.80 12.00 157.46 12.66 ;
      LAYER Metal6 ;
        RECT 156.80 12.00 157.46 12.66 ;
      LAYER Metal3 ;
        RECT 156.80 12.00 157.46 12.66 ;
      LAYER Metal4 ;
        RECT 156.80 12.00 157.46 12.66 ;
    END
  END Q[13]
  PIN Q[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 175.20 12.00 175.86 12.66 ;
      LAYER Metal6 ;
        RECT 175.20 12.00 175.86 12.66 ;
      LAYER Metal3 ;
        RECT 175.20 12.00 175.86 12.66 ;
      LAYER Metal4 ;
        RECT 175.20 12.00 175.86 12.66 ;
    END
  END Q[14]
  PIN Q[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 178.08 12.00 178.74 12.66 ;
      LAYER Metal6 ;
        RECT 178.08 12.00 178.74 12.66 ;
      LAYER Metal3 ;
        RECT 178.08 12.00 178.74 12.66 ;
      LAYER Metal4 ;
        RECT 178.08 12.00 178.74 12.66 ;
    END
  END Q[15]
  PIN Q[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 248.22 12.00 248.88 12.66 ;
      LAYER Metal6 ;
        RECT 248.22 12.00 248.88 12.66 ;
      LAYER Metal3 ;
        RECT 248.22 12.00 248.88 12.66 ;
      LAYER Metal4 ;
        RECT 248.22 12.00 248.88 12.66 ;
    END
  END Q[16]
  PIN Q[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 251.10 12.00 251.76 12.66 ;
      LAYER Metal6 ;
        RECT 251.10 12.00 251.76 12.66 ;
      LAYER Metal3 ;
        RECT 251.10 12.00 251.76 12.66 ;
      LAYER Metal4 ;
        RECT 251.10 12.00 251.76 12.66 ;
    END
  END Q[17]
  PIN Q[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 269.50 12.00 270.17 12.66 ;
      LAYER Metal6 ;
        RECT 269.50 12.00 270.17 12.66 ;
      LAYER Metal3 ;
        RECT 269.50 12.00 270.17 12.66 ;
      LAYER Metal4 ;
        RECT 269.50 12.00 270.17 12.66 ;
    END
  END Q[18]
  PIN Q[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 272.38 12.00 273.05 12.66 ;
      LAYER Metal6 ;
        RECT 272.38 12.00 273.05 12.66 ;
      LAYER Metal3 ;
        RECT 272.38 12.00 273.05 12.66 ;
      LAYER Metal4 ;
        RECT 272.38 12.00 273.05 12.66 ;
    END
  END Q[19]
  PIN Q[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 25.94 12.00 26.60 12.66 ;
      LAYER Metal6 ;
        RECT 25.94 12.00 26.60 12.66 ;
      LAYER Metal3 ;
        RECT 25.94 12.00 26.60 12.66 ;
      LAYER Metal4 ;
        RECT 25.94 12.00 26.60 12.66 ;
    END
  END Q[1]
  PIN Q[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 291.85 12.00 292.50 12.66 ;
      LAYER Metal6 ;
        RECT 291.85 12.00 292.50 12.66 ;
      LAYER Metal3 ;
        RECT 291.85 12.00 292.50 12.66 ;
      LAYER Metal4 ;
        RECT 291.85 12.00 292.50 12.66 ;
    END
  END Q[20]
  PIN Q[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 294.73 12.00 295.38 12.66 ;
      LAYER Metal6 ;
        RECT 294.73 12.00 295.38 12.66 ;
      LAYER Metal3 ;
        RECT 294.73 12.00 295.38 12.66 ;
      LAYER Metal4 ;
        RECT 294.73 12.00 295.38 12.66 ;
    END
  END Q[21]
  PIN Q[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 313.12 12.00 313.79 12.66 ;
      LAYER Metal6 ;
        RECT 313.12 12.00 313.79 12.66 ;
      LAYER Metal3 ;
        RECT 313.12 12.00 313.79 12.66 ;
      LAYER Metal4 ;
        RECT 313.12 12.00 313.79 12.66 ;
    END
  END Q[22]
  PIN Q[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 316.00 12.00 316.67 12.66 ;
      LAYER Metal6 ;
        RECT 316.00 12.00 316.67 12.66 ;
      LAYER Metal3 ;
        RECT 316.00 12.00 316.67 12.66 ;
      LAYER Metal4 ;
        RECT 316.00 12.00 316.67 12.66 ;
    END
  END Q[23]
  PIN Q[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 335.46 12.00 336.12 12.66 ;
      LAYER Metal6 ;
        RECT 335.46 12.00 336.12 12.66 ;
      LAYER Metal3 ;
        RECT 335.46 12.00 336.12 12.66 ;
      LAYER Metal4 ;
        RECT 335.46 12.00 336.12 12.66 ;
    END
  END Q[24]
  PIN Q[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 338.35 12.00 339.00 12.66 ;
      LAYER Metal6 ;
        RECT 338.35 12.00 339.00 12.66 ;
      LAYER Metal3 ;
        RECT 338.35 12.00 339.00 12.66 ;
      LAYER Metal4 ;
        RECT 338.35 12.00 339.00 12.66 ;
    END
  END Q[25]
  PIN Q[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 356.75 12.00 357.40 12.66 ;
      LAYER Metal6 ;
        RECT 356.75 12.00 357.40 12.66 ;
      LAYER Metal3 ;
        RECT 356.75 12.00 357.40 12.66 ;
      LAYER Metal4 ;
        RECT 356.75 12.00 357.40 12.66 ;
    END
  END Q[26]
  PIN Q[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 359.62 12.00 360.29 12.66 ;
      LAYER Metal6 ;
        RECT 359.62 12.00 360.29 12.66 ;
      LAYER Metal3 ;
        RECT 359.62 12.00 360.29 12.66 ;
      LAYER Metal4 ;
        RECT 359.62 12.00 360.29 12.66 ;
    END
  END Q[27]
  PIN Q[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 379.08 12.00 379.75 12.66 ;
      LAYER Metal6 ;
        RECT 379.08 12.00 379.75 12.66 ;
      LAYER Metal3 ;
        RECT 379.08 12.00 379.75 12.66 ;
      LAYER Metal4 ;
        RECT 379.08 12.00 379.75 12.66 ;
    END
  END Q[28]
  PIN Q[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 381.96 12.00 382.62 12.66 ;
      LAYER Metal6 ;
        RECT 381.96 12.00 382.62 12.66 ;
      LAYER Metal3 ;
        RECT 381.96 12.00 382.62 12.66 ;
      LAYER Metal4 ;
        RECT 381.96 12.00 382.62 12.66 ;
    END
  END Q[29]
  PIN Q[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 44.34 12.00 45.00 12.66 ;
      LAYER Metal6 ;
        RECT 44.34 12.00 45.00 12.66 ;
      LAYER Metal3 ;
        RECT 44.34 12.00 45.00 12.66 ;
      LAYER Metal4 ;
        RECT 44.34 12.00 45.00 12.66 ;
    END
  END Q[2]
  PIN Q[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 400.37 12.00 401.02 12.66 ;
      LAYER Metal6 ;
        RECT 400.37 12.00 401.02 12.66 ;
      LAYER Metal3 ;
        RECT 400.37 12.00 401.02 12.66 ;
      LAYER Metal4 ;
        RECT 400.37 12.00 401.02 12.66 ;
    END
  END Q[30]
  PIN Q[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 403.25 12.00 403.90 12.66 ;
      LAYER Metal6 ;
        RECT 403.25 12.00 403.90 12.66 ;
      LAYER Metal3 ;
        RECT 403.25 12.00 403.90 12.66 ;
      LAYER Metal4 ;
        RECT 403.25 12.00 403.90 12.66 ;
    END
  END Q[31]
  PIN Q[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 47.22 12.00 47.88 12.66 ;
      LAYER Metal6 ;
        RECT 47.22 12.00 47.88 12.66 ;
      LAYER Metal3 ;
        RECT 47.22 12.00 47.88 12.66 ;
      LAYER Metal4 ;
        RECT 47.22 12.00 47.88 12.66 ;
    END
  END Q[3]
  PIN Q[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 66.68 12.00 67.34 12.66 ;
      LAYER Metal6 ;
        RECT 66.68 12.00 67.34 12.66 ;
      LAYER Metal3 ;
        RECT 66.68 12.00 67.34 12.66 ;
      LAYER Metal4 ;
        RECT 66.68 12.00 67.34 12.66 ;
    END
  END Q[4]
  PIN Q[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 69.56 12.00 70.22 12.66 ;
      LAYER Metal6 ;
        RECT 69.56 12.00 70.22 12.66 ;
      LAYER Metal3 ;
        RECT 69.56 12.00 70.22 12.66 ;
      LAYER Metal4 ;
        RECT 69.56 12.00 70.22 12.66 ;
    END
  END Q[5]
  PIN Q[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 87.96 12.00 88.62 12.66 ;
      LAYER Metal6 ;
        RECT 87.96 12.00 88.62 12.66 ;
      LAYER Metal3 ;
        RECT 87.96 12.00 88.62 12.66 ;
      LAYER Metal4 ;
        RECT 87.96 12.00 88.62 12.66 ;
    END
  END Q[6]
  PIN Q[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 90.84 12.00 91.50 12.66 ;
      LAYER Metal6 ;
        RECT 90.84 12.00 91.50 12.66 ;
      LAYER Metal3 ;
        RECT 90.84 12.00 91.50 12.66 ;
      LAYER Metal4 ;
        RECT 90.84 12.00 91.50 12.66 ;
    END
  END Q[7]
  PIN Q[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 110.30 12.00 110.96 12.66 ;
      LAYER Metal6 ;
        RECT 110.30 12.00 110.96 12.66 ;
      LAYER Metal3 ;
        RECT 110.30 12.00 110.96 12.66 ;
      LAYER Metal4 ;
        RECT 110.30 12.00 110.96 12.66 ;
    END
  END Q[8]
  PIN Q[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 113.18 12.00 113.84 12.66 ;
      LAYER Metal6 ;
        RECT 113.18 12.00 113.84 12.66 ;
      LAYER Metal3 ;
        RECT 113.18 12.00 113.84 12.66 ;
      LAYER Metal4 ;
        RECT 113.18 12.00 113.84 12.66 ;
    END
  END Q[9]
  PIN WE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 234.48 12.00 235.14 12.66 ;
      LAYER Metal6 ;
        RECT 234.48 12.00 235.14 12.66 ;
      LAYER Metal3 ;
        RECT 234.48 12.00 235.14 12.66 ;
      LAYER Metal4 ;
        RECT 234.48 12.00 235.14 12.66 ;
    END
  END WE
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE RING ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 109.22 426.96 114.22 ;
        RECT 0.00 0.00 426.96 5.00 ;
      LAYER Metal2 ;
        RECT 421.96 0.00 426.96 114.22 ;
        RECT 0.00 0.00 5.00 114.22 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE RING ;
    PORT
      LAYER Metal1 ;
        RECT 5.60 103.61 421.37 108.61 ;
        RECT 5.60 5.60 421.37 10.60 ;
      LAYER Metal2 ;
        RECT 416.37 5.60 421.37 108.61 ;
        RECT 5.60 5.60 10.60 108.61 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      RECT 12.00 12.00 415.01 102.02 ;
    LAYER Metal2 ;
      RECT 12.00 12.00 415.01 102.02 ;
    LAYER Metal3 ;
#      RECT 12.00 12.00 415.01 102.02 ;
        RECT 12.84 12.84 415.01 102.02 ;
        RECT 12.00 12.00 20.30 46.86 ;
        RECT 21.32 12.00 22.88 102.02 ;
        RECT 23.90 12.00 25.76 102.02 ;
        RECT 26.78 12.00 28.34 102.02 ;
        RECT 29.36 12.00 41.58 102.02 ;
        RECT 42.60 12.00 44.16 102.02 ;
        RECT 45.18 12.00 47.04 102.02 ;
        RECT 48.06 12.00 49.62 102.02 ;
        RECT 50.64 12.00 63.92 102.02 ;
        RECT 64.94 12.00 66.50 102.02 ;
        RECT 67.52 12.00 69.38 102.02 ;
        RECT 70.40 12.00 71.96 102.02 ;
        RECT 72.98 12.00 85.20 102.02 ;
        RECT 86.22 12.00 87.78 102.02 ;
        RECT 88.80 12.00 90.66 102.02 ;
        RECT 91.68 12.00 93.24 102.02 ;
        RECT 94.26 12.00 107.54 102.02 ;
        RECT 108.56 12.00 110.12 102.02 ;
        RECT 111.14 12.00 113.00 102.02 ;
        RECT 114.02 12.00 115.58 102.02 ;
        RECT 116.60 12.00 128.82 102.02 ;
        RECT 129.84 12.00 131.40 102.02 ;
        RECT 132.42 12.00 134.28 102.02 ;
        RECT 135.30 12.00 136.86 102.02 ;
        RECT 137.88 12.00 151.16 102.02 ;
        RECT 152.18 12.00 153.74 102.02 ;
        RECT 154.76 12.00 156.62 102.02 ;
        RECT 157.64 12.00 159.20 102.02 ;
        RECT 160.22 12.00 172.44 102.02 ;
        RECT 173.46 12.00 175.02 102.02 ;
        RECT 176.04 12.00 177.90 102.02 ;
        RECT 178.92 12.00 180.48 102.02 ;
        RECT 181.50 12.00 228.26 102.02 ;
        RECT 229.27 12.00 234.30 102.02 ;
        RECT 235.32 12.00 238.00 102.02 ;
        RECT 239.02 12.00 245.47 102.02 ;
        RECT 246.49 12.00 248.04 102.02 ;
        RECT 249.06 12.00 250.92 102.02 ;
        RECT 251.94 12.00 253.51 102.02 ;
        RECT 254.52 12.00 266.75 102.02 ;
        RECT 267.76 12.00 269.32 102.02 ;
        RECT 270.35 12.00 272.20 102.02 ;
        RECT 273.23 12.00 274.78 102.02 ;
        RECT 275.80 12.00 289.08 102.02 ;
        RECT 290.11 12.00 291.67 102.02 ;
        RECT 292.68 12.00 294.55 102.02 ;
        RECT 295.56 12.00 297.13 102.02 ;
        RECT 298.14 12.00 310.37 102.02 ;
        RECT 311.38 12.00 312.94 102.02 ;
        RECT 313.97 12.00 315.82 102.02 ;
        RECT 316.85 12.00 318.40 102.02 ;
        RECT 319.43 12.00 332.70 102.02 ;
        RECT 333.73 12.00 335.28 102.02 ;
        RECT 336.30 12.00 338.17 102.02 ;
        RECT 339.18 12.00 340.75 102.02 ;
        RECT 341.76 12.00 353.99 102.02 ;
        RECT 355.00 12.00 356.57 102.02 ;
        RECT 357.58 12.00 359.44 102.02 ;
        RECT 360.47 12.00 362.02 102.02 ;
        RECT 363.05 12.00 376.32 102.02 ;
        RECT 377.35 12.00 378.90 102.02 ;
        RECT 379.93 12.00 381.78 102.02 ;
        RECT 382.80 12.00 384.37 102.02 ;
        RECT 385.38 12.00 397.61 102.02 ;
        RECT 398.62 12.00 400.19 102.02 ;
        RECT 401.20 12.00 403.07 102.02 ;
        RECT 404.08 12.00 405.64 102.02 ;
        RECT 406.67 12.00 415.01 102.02 ;
        RECT 12.00 47.88 415.01 49.88 ;
        RECT 12.00 50.90 415.01 56.00 ;
        RECT 12.00 57.02 415.01 59.10 ;
        RECT 12.00 60.12 415.01 62.12 ;
        RECT 12.00 63.14 415.01 68.24 ;
        RECT 12.00 69.26 415.01 71.34 ;
        RECT 12.00 72.36 415.01 77.46 ;
        RECT 12.00 78.48 415.01 102.02 ;
    LAYER Metal4 ;
#      RECT 12.00 12.00 415.01 102.02 ;
        RECT 12.84 12.84 415.01 102.02 ;
        RECT 12.00 12.00 20.30 46.86 ;
        RECT 21.32 12.00 22.88 102.02 ;
        RECT 23.90 12.00 25.76 102.02 ;
        RECT 26.78 12.00 28.34 102.02 ;
        RECT 29.36 12.00 41.58 102.02 ;
        RECT 42.60 12.00 44.16 102.02 ;
        RECT 45.18 12.00 47.04 102.02 ;
        RECT 48.06 12.00 49.62 102.02 ;
        RECT 50.64 12.00 63.92 102.02 ;
        RECT 64.94 12.00 66.50 102.02 ;
        RECT 67.52 12.00 69.38 102.02 ;
        RECT 70.40 12.00 71.96 102.02 ;
        RECT 72.98 12.00 85.20 102.02 ;
        RECT 86.22 12.00 87.78 102.02 ;
        RECT 88.80 12.00 90.66 102.02 ;
        RECT 91.68 12.00 93.24 102.02 ;
        RECT 94.26 12.00 107.54 102.02 ;
        RECT 108.56 12.00 110.12 102.02 ;
        RECT 111.14 12.00 113.00 102.02 ;
        RECT 114.02 12.00 115.58 102.02 ;
        RECT 116.60 12.00 128.82 102.02 ;
        RECT 129.84 12.00 131.40 102.02 ;
        RECT 132.42 12.00 134.28 102.02 ;
        RECT 135.30 12.00 136.86 102.02 ;
        RECT 137.88 12.00 151.16 102.02 ;
        RECT 152.18 12.00 153.74 102.02 ;
        RECT 154.76 12.00 156.62 102.02 ;
        RECT 157.64 12.00 159.20 102.02 ;
        RECT 160.22 12.00 172.44 102.02 ;
        RECT 173.46 12.00 175.02 102.02 ;
        RECT 176.04 12.00 177.90 102.02 ;
        RECT 178.92 12.00 180.48 102.02 ;
        RECT 181.50 12.00 228.26 102.02 ;
        RECT 229.27 12.00 234.30 102.02 ;
        RECT 235.32 12.00 238.00 102.02 ;
        RECT 239.02 12.00 245.47 102.02 ;
        RECT 246.49 12.00 248.04 102.02 ;
        RECT 249.06 12.00 250.92 102.02 ;
        RECT 251.94 12.00 253.51 102.02 ;
        RECT 254.52 12.00 266.75 102.02 ;
        RECT 267.76 12.00 269.32 102.02 ;
        RECT 270.35 12.00 272.20 102.02 ;
        RECT 273.23 12.00 274.78 102.02 ;
        RECT 275.80 12.00 289.08 102.02 ;
        RECT 290.11 12.00 291.67 102.02 ;
        RECT 292.68 12.00 294.55 102.02 ;
        RECT 295.56 12.00 297.13 102.02 ;
        RECT 298.14 12.00 310.37 102.02 ;
        RECT 311.38 12.00 312.94 102.02 ;
        RECT 313.97 12.00 315.82 102.02 ;
        RECT 316.85 12.00 318.40 102.02 ;
        RECT 319.43 12.00 332.70 102.02 ;
        RECT 333.73 12.00 335.28 102.02 ;
        RECT 336.30 12.00 338.17 102.02 ;
        RECT 339.18 12.00 340.75 102.02 ;
        RECT 341.76 12.00 353.99 102.02 ;
        RECT 355.00 12.00 356.57 102.02 ;
        RECT 357.58 12.00 359.44 102.02 ;
        RECT 360.47 12.00 362.02 102.02 ;
        RECT 363.05 12.00 376.32 102.02 ;
        RECT 377.35 12.00 378.90 102.02 ;
        RECT 379.93 12.00 381.78 102.02 ;
        RECT 382.80 12.00 384.37 102.02 ;
        RECT 385.38 12.00 397.61 102.02 ;
        RECT 398.62 12.00 400.19 102.02 ;
        RECT 401.20 12.00 403.07 102.02 ;
        RECT 404.08 12.00 405.64 102.02 ;
        RECT 406.67 12.00 415.01 102.02 ;
        RECT 12.00 47.88 415.01 49.88 ;
        RECT 12.00 50.90 415.01 56.00 ;
        RECT 12.00 57.02 415.01 59.10 ;
        RECT 12.00 60.12 415.01 62.12 ;
        RECT 12.00 63.14 415.01 68.24 ;
        RECT 12.00 69.26 415.01 71.34 ;
        RECT 12.00 72.36 415.01 77.46 ;
        RECT 12.00 78.48 415.01 102.02 ;
    LAYER Metal5 ;
#      RECT 12.00 12.00 415.01 102.02 ;
        RECT 12.84 12.84 415.01 102.02 ;
        RECT 12.00 12.00 20.30 46.86 ;
        RECT 21.32 12.00 22.88 102.02 ;
        RECT 23.90 12.00 25.76 102.02 ;
        RECT 26.78 12.00 28.34 102.02 ;
        RECT 29.36 12.00 41.58 102.02 ;
        RECT 42.60 12.00 44.16 102.02 ;
        RECT 45.18 12.00 47.04 102.02 ;
        RECT 48.06 12.00 49.62 102.02 ;
        RECT 50.64 12.00 63.92 102.02 ;
        RECT 64.94 12.00 66.50 102.02 ;
        RECT 67.52 12.00 69.38 102.02 ;
        RECT 70.40 12.00 71.96 102.02 ;
        RECT 72.98 12.00 85.20 102.02 ;
        RECT 86.22 12.00 87.78 102.02 ;
        RECT 88.80 12.00 90.66 102.02 ;
        RECT 91.68 12.00 93.24 102.02 ;
        RECT 94.26 12.00 107.54 102.02 ;
        RECT 108.56 12.00 110.12 102.02 ;
        RECT 111.14 12.00 113.00 102.02 ;
        RECT 114.02 12.00 115.58 102.02 ;
        RECT 116.60 12.00 128.82 102.02 ;
        RECT 129.84 12.00 131.40 102.02 ;
        RECT 132.42 12.00 134.28 102.02 ;
        RECT 135.30 12.00 136.86 102.02 ;
        RECT 137.88 12.00 151.16 102.02 ;
        RECT 152.18 12.00 153.74 102.02 ;
        RECT 154.76 12.00 156.62 102.02 ;
        RECT 157.64 12.00 159.20 102.02 ;
        RECT 160.22 12.00 172.44 102.02 ;
        RECT 173.46 12.00 175.02 102.02 ;
        RECT 176.04 12.00 177.90 102.02 ;
        RECT 178.92 12.00 180.48 102.02 ;
        RECT 181.50 12.00 228.26 102.02 ;
        RECT 229.27 12.00 234.30 102.02 ;
        RECT 235.32 12.00 238.00 102.02 ;
        RECT 239.02 12.00 245.47 102.02 ;
        RECT 246.49 12.00 248.04 102.02 ;
        RECT 249.06 12.00 250.92 102.02 ;
        RECT 251.94 12.00 253.51 102.02 ;
        RECT 254.52 12.00 266.75 102.02 ;
        RECT 267.76 12.00 269.32 102.02 ;
        RECT 270.35 12.00 272.20 102.02 ;
        RECT 273.23 12.00 274.78 102.02 ;
        RECT 275.80 12.00 289.08 102.02 ;
        RECT 290.11 12.00 291.67 102.02 ;
        RECT 292.68 12.00 294.55 102.02 ;
        RECT 295.56 12.00 297.13 102.02 ;
        RECT 298.14 12.00 310.37 102.02 ;
        RECT 311.38 12.00 312.94 102.02 ;
        RECT 313.97 12.00 315.82 102.02 ;
        RECT 316.85 12.00 318.40 102.02 ;
        RECT 319.43 12.00 332.70 102.02 ;
        RECT 333.73 12.00 335.28 102.02 ;
        RECT 336.30 12.00 338.17 102.02 ;
        RECT 339.18 12.00 340.75 102.02 ;
        RECT 341.76 12.00 353.99 102.02 ;
        RECT 355.00 12.00 356.57 102.02 ;
        RECT 357.58 12.00 359.44 102.02 ;
        RECT 360.47 12.00 362.02 102.02 ;
        RECT 363.05 12.00 376.32 102.02 ;
        RECT 377.35 12.00 378.90 102.02 ;
        RECT 379.93 12.00 381.78 102.02 ;
        RECT 382.80 12.00 384.37 102.02 ;
        RECT 385.38 12.00 397.61 102.02 ;
        RECT 398.62 12.00 400.19 102.02 ;
        RECT 401.20 12.00 403.07 102.02 ;
        RECT 404.08 12.00 405.64 102.02 ;
        RECT 406.67 12.00 415.01 102.02 ;
        RECT 12.00 47.88 415.01 49.88 ;
        RECT 12.00 50.90 415.01 56.00 ;
        RECT 12.00 57.02 415.01 59.10 ;
        RECT 12.00 60.12 415.01 62.12 ;
        RECT 12.00 63.14 415.01 68.24 ;
        RECT 12.00 69.26 415.01 71.34 ;
        RECT 12.00 72.36 415.01 77.46 ;
        RECT 12.00 78.48 415.01 102.02 ;
    LAYER Metal6 ;
#      RECT 12.00 12.00 415.01 102.02 ;
        RECT 12.84 12.84 415.01 102.02 ;
        RECT 12.00 12.00 20.30 46.86 ;
        RECT 21.32 12.00 22.88 102.02 ;
        RECT 23.90 12.00 25.76 102.02 ;
        RECT 26.78 12.00 28.34 102.02 ;
        RECT 29.36 12.00 41.58 102.02 ;
        RECT 42.60 12.00 44.16 102.02 ;
        RECT 45.18 12.00 47.04 102.02 ;
        RECT 48.06 12.00 49.62 102.02 ;
        RECT 50.64 12.00 63.92 102.02 ;
        RECT 64.94 12.00 66.50 102.02 ;
        RECT 67.52 12.00 69.38 102.02 ;
        RECT 70.40 12.00 71.96 102.02 ;
        RECT 72.98 12.00 85.20 102.02 ;
        RECT 86.22 12.00 87.78 102.02 ;
        RECT 88.80 12.00 90.66 102.02 ;
        RECT 91.68 12.00 93.24 102.02 ;
        RECT 94.26 12.00 107.54 102.02 ;
        RECT 108.56 12.00 110.12 102.02 ;
        RECT 111.14 12.00 113.00 102.02 ;
        RECT 114.02 12.00 115.58 102.02 ;
        RECT 116.60 12.00 128.82 102.02 ;
        RECT 129.84 12.00 131.40 102.02 ;
        RECT 132.42 12.00 134.28 102.02 ;
        RECT 135.30 12.00 136.86 102.02 ;
        RECT 137.88 12.00 151.16 102.02 ;
        RECT 152.18 12.00 153.74 102.02 ;
        RECT 154.76 12.00 156.62 102.02 ;
        RECT 157.64 12.00 159.20 102.02 ;
        RECT 160.22 12.00 172.44 102.02 ;
        RECT 173.46 12.00 175.02 102.02 ;
        RECT 176.04 12.00 177.90 102.02 ;
        RECT 178.92 12.00 180.48 102.02 ;
        RECT 181.50 12.00 228.26 102.02 ;
        RECT 229.27 12.00 234.30 102.02 ;
        RECT 235.32 12.00 238.00 102.02 ;
        RECT 239.02 12.00 245.47 102.02 ;
        RECT 246.49 12.00 248.04 102.02 ;
        RECT 249.06 12.00 250.92 102.02 ;
        RECT 251.94 12.00 253.51 102.02 ;
        RECT 254.52 12.00 266.75 102.02 ;
        RECT 267.76 12.00 269.32 102.02 ;
        RECT 270.35 12.00 272.20 102.02 ;
        RECT 273.23 12.00 274.78 102.02 ;
        RECT 275.80 12.00 289.08 102.02 ;
        RECT 290.11 12.00 291.67 102.02 ;
        RECT 292.68 12.00 294.55 102.02 ;
        RECT 295.56 12.00 297.13 102.02 ;
        RECT 298.14 12.00 310.37 102.02 ;
        RECT 311.38 12.00 312.94 102.02 ;
        RECT 313.97 12.00 315.82 102.02 ;
        RECT 316.85 12.00 318.40 102.02 ;
        RECT 319.43 12.00 332.70 102.02 ;
        RECT 333.73 12.00 335.28 102.02 ;
        RECT 336.30 12.00 338.17 102.02 ;
        RECT 339.18 12.00 340.75 102.02 ;
        RECT 341.76 12.00 353.99 102.02 ;
        RECT 355.00 12.00 356.57 102.02 ;
        RECT 357.58 12.00 359.44 102.02 ;
        RECT 360.47 12.00 362.02 102.02 ;
        RECT 363.05 12.00 376.32 102.02 ;
        RECT 377.35 12.00 378.90 102.02 ;
        RECT 379.93 12.00 381.78 102.02 ;
        RECT 382.80 12.00 384.37 102.02 ;
        RECT 385.38 12.00 397.61 102.02 ;
        RECT 398.62 12.00 400.19 102.02 ;
        RECT 401.20 12.00 403.07 102.02 ;
        RECT 404.08 12.00 405.64 102.02 ;
        RECT 406.67 12.00 415.01 102.02 ;
        RECT 12.00 47.88 415.01 49.88 ;
        RECT 12.00 50.90 415.01 56.00 ;
        RECT 12.00 57.02 415.01 59.10 ;
        RECT 12.00 60.12 415.01 62.12 ;
        RECT 12.00 63.14 415.01 68.24 ;
        RECT 12.00 69.26 415.01 71.34 ;
        RECT 12.00 72.36 415.01 77.46 ;
        RECT 12.00 78.48 415.01 102.02 ;
  END
END MEM1

MACRO MEM2
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN MEM2 0 0 ;
  SIZE 423.015 BY 145.035 ;
  SYMMETRY X Y R90 ;
  PIN A1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12.00 102.42 12.66 103.08 ;
      LAYER Metal6 ;
        RECT 12.00 102.42 12.66 103.08 ;
      LAYER Metal3 ;
        RECT 12.00 102.42 12.66 103.08 ;
      LAYER Metal4 ;
        RECT 12.00 102.42 12.66 103.08 ;
    END
  END A1[0]
  PIN A1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12.00 96.30 12.66 96.96 ;
      LAYER Metal6 ;
        RECT 12.00 96.30 12.66 96.96 ;
      LAYER Metal3 ;
        RECT 12.00 96.30 12.66 96.96 ;
      LAYER Metal4 ;
        RECT 12.00 96.30 12.66 96.96 ;
    END
  END A1[1]
  PIN A1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12.00 87.08 12.66 87.74 ;
      LAYER Metal6 ;
        RECT 12.00 87.08 12.66 87.74 ;
      LAYER Metal3 ;
        RECT 12.00 87.08 12.66 87.74 ;
      LAYER Metal4 ;
        RECT 12.00 87.08 12.66 87.74 ;
    END
  END A1[2]
  PIN A1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12.00 84.06 12.66 84.72 ;
      LAYER Metal6 ;
        RECT 12.00 84.06 12.66 84.72 ;
      LAYER Metal3 ;
        RECT 12.00 84.06 12.66 84.72 ;
      LAYER Metal4 ;
        RECT 12.00 84.06 12.66 84.72 ;
    END
  END A1[3]
  PIN A1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12.00 80.96 12.66 81.62 ;
      LAYER Metal6 ;
        RECT 12.00 80.96 12.66 81.62 ;
      LAYER Metal3 ;
        RECT 12.00 80.96 12.66 81.62 ;
      LAYER Metal4 ;
        RECT 12.00 80.96 12.66 81.62 ;
    END
  END A1[4]
  PIN A1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12.00 74.84 12.66 75.50 ;
      LAYER Metal6 ;
        RECT 12.00 74.84 12.66 75.50 ;
      LAYER Metal3 ;
        RECT 12.00 74.84 12.66 75.50 ;
      LAYER Metal4 ;
        RECT 12.00 74.84 12.66 75.50 ;
    END
  END A1[5]
  PIN A1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12.00 71.82 12.66 72.48 ;
      LAYER Metal6 ;
        RECT 12.00 71.82 12.66 72.48 ;
      LAYER Metal3 ;
        RECT 12.00 71.82 12.66 72.48 ;
      LAYER Metal4 ;
        RECT 12.00 71.82 12.66 72.48 ;
    END
  END A1[6]
  PIN A2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12.00 36.40 12.66 37.06 ;
      LAYER Metal6 ;
        RECT 12.00 36.40 12.66 37.06 ;
      LAYER Metal3 ;
        RECT 12.00 36.40 12.66 37.06 ;
      LAYER Metal4 ;
        RECT 12.00 36.40 12.66 37.06 ;
    END
  END A2[0]
  PIN A2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12.00 42.52 12.66 43.18 ;
      LAYER Metal6 ;
        RECT 12.00 42.52 12.66 43.18 ;
      LAYER Metal3 ;
        RECT 12.00 42.52 12.66 43.18 ;
      LAYER Metal4 ;
        RECT 12.00 42.52 12.66 43.18 ;
    END
  END A2[1]
  PIN A2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12.00 51.74 12.66 52.40 ;
      LAYER Metal6 ;
        RECT 12.00 51.74 12.66 52.40 ;
      LAYER Metal3 ;
        RECT 12.00 51.74 12.66 52.40 ;
      LAYER Metal4 ;
        RECT 12.00 51.74 12.66 52.40 ;
    END
  END A2[2]
  PIN A2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12.00 54.76 12.66 55.42 ;
      LAYER Metal6 ;
        RECT 12.00 54.76 12.66 55.42 ;
      LAYER Metal3 ;
        RECT 12.00 54.76 12.66 55.42 ;
      LAYER Metal4 ;
        RECT 12.00 54.76 12.66 55.42 ;
    END
  END A2[3]
  PIN A2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12.00 57.86 12.66 58.52 ;
      LAYER Metal6 ;
        RECT 12.00 57.86 12.66 58.52 ;
      LAYER Metal3 ;
        RECT 12.00 57.86 12.66 58.52 ;
      LAYER Metal4 ;
        RECT 12.00 57.86 12.66 58.52 ;
    END
  END A2[4]
  PIN A2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12.00 63.98 12.66 64.64 ;
      LAYER Metal6 ;
        RECT 12.00 63.98 12.66 64.64 ;
      LAYER Metal3 ;
        RECT 12.00 63.98 12.66 64.64 ;
      LAYER Metal4 ;
        RECT 12.00 63.98 12.66 64.64 ;
    END
  END A2[5]
  PIN A2[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12.00 67.00 12.66 67.66 ;
      LAYER Metal6 ;
        RECT 12.00 67.00 12.66 67.66 ;
      LAYER Metal3 ;
        RECT 12.00 67.00 12.66 67.66 ;
      LAYER Metal4 ;
        RECT 12.00 67.00 12.66 67.66 ;
    END
  END A2[6]
  PIN CE1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 210.28 12.00 210.94 12.66 ;
      LAYER Metal6 ;
        RECT 210.28 12.00 210.94 12.66 ;
      LAYER Metal3 ;
        RECT 210.28 12.00 210.94 12.66 ;
      LAYER Metal4 ;
        RECT 210.28 12.00 210.94 12.66 ;
    END
  END CE1
  PIN CE2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 196.36 12.00 197.02 12.66 ;
      LAYER Metal6 ;
        RECT 196.36 12.00 197.02 12.66 ;
      LAYER Metal3 ;
        RECT 196.36 12.00 197.02 12.66 ;
      LAYER Metal4 ;
        RECT 196.36 12.00 197.02 12.66 ;
    END
  END CE2
  PIN CK1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 218.91 12.00 219.56 12.66 ;
      LAYER Metal6 ;
        RECT 218.91 12.00 219.56 12.66 ;
      LAYER Metal3 ;
        RECT 218.91 12.00 219.56 12.66 ;
      LAYER Metal4 ;
        RECT 218.91 12.00 219.56 12.66 ;
    END
  END CK1
  PIN CK2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 187.74 12.00 188.40 12.66 ;
      LAYER Metal6 ;
        RECT 187.74 12.00 188.40 12.66 ;
      LAYER Metal3 ;
        RECT 187.74 12.00 188.40 12.66 ;
      LAYER Metal4 ;
        RECT 187.74 12.00 188.40 12.66 ;
    END
  END CK2
  PIN D1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 15.86 12.00 16.52 12.66 ;
      LAYER Metal6 ;
        RECT 15.86 12.00 16.52 12.66 ;
      LAYER Metal3 ;
        RECT 15.86 12.00 16.52 12.66 ;
      LAYER Metal4 ;
        RECT 15.86 12.00 16.52 12.66 ;
    END
  END D1[0]
  PIN D1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 122.26 12.00 122.92 12.66 ;
      LAYER Metal6 ;
        RECT 122.26 12.00 122.92 12.66 ;
      LAYER Metal3 ;
        RECT 122.26 12.00 122.92 12.66 ;
      LAYER Metal4 ;
        RECT 122.26 12.00 122.92 12.66 ;
    END
  END D1[10]
  PIN D1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 142.40 12.00 143.06 12.66 ;
      LAYER Metal6 ;
        RECT 142.40 12.00 143.06 12.66 ;
      LAYER Metal3 ;
        RECT 142.40 12.00 143.06 12.66 ;
      LAYER Metal4 ;
        RECT 142.40 12.00 143.06 12.66 ;
    END
  END D1[11]
  PIN D1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 143.54 12.00 144.20 12.66 ;
      LAYER Metal6 ;
        RECT 143.54 12.00 144.20 12.66 ;
      LAYER Metal3 ;
        RECT 143.54 12.00 144.20 12.66 ;
      LAYER Metal4 ;
        RECT 143.54 12.00 144.20 12.66 ;
    END
  END D1[12]
  PIN D1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 163.68 12.00 164.34 12.66 ;
      LAYER Metal6 ;
        RECT 163.68 12.00 164.34 12.66 ;
      LAYER Metal3 ;
        RECT 163.68 12.00 164.34 12.66 ;
      LAYER Metal4 ;
        RECT 163.68 12.00 164.34 12.66 ;
    END
  END D1[13]
  PIN D1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 164.82 12.00 165.48 12.66 ;
      LAYER Metal6 ;
        RECT 164.82 12.00 165.48 12.66 ;
      LAYER Metal3 ;
        RECT 164.82 12.00 165.48 12.66 ;
      LAYER Metal4 ;
        RECT 164.82 12.00 165.48 12.66 ;
    END
  END D1[14]
  PIN D1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 184.96 12.00 185.62 12.66 ;
      LAYER Metal6 ;
        RECT 184.96 12.00 185.62 12.66 ;
      LAYER Metal3 ;
        RECT 184.96 12.00 185.62 12.66 ;
      LAYER Metal4 ;
        RECT 184.96 12.00 185.62 12.66 ;
    END
  END D1[15]
  PIN D1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 221.68 12.00 222.34 12.66 ;
      LAYER Metal6 ;
        RECT 221.68 12.00 222.34 12.66 ;
      LAYER Metal3 ;
        RECT 221.68 12.00 222.34 12.66 ;
      LAYER Metal4 ;
        RECT 221.68 12.00 222.34 12.66 ;
    END
  END D1[16]
  PIN D1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 241.82 12.00 242.48 12.66 ;
      LAYER Metal6 ;
        RECT 241.82 12.00 242.48 12.66 ;
      LAYER Metal3 ;
        RECT 241.82 12.00 242.48 12.66 ;
      LAYER Metal4 ;
        RECT 241.82 12.00 242.48 12.66 ;
    END
  END D1[17]
  PIN D1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 242.96 12.00 243.62 12.66 ;
      LAYER Metal6 ;
        RECT 242.96 12.00 243.62 12.66 ;
      LAYER Metal3 ;
        RECT 242.96 12.00 243.62 12.66 ;
      LAYER Metal4 ;
        RECT 242.96 12.00 243.62 12.66 ;
    END
  END D1[18]
  PIN D1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 263.10 12.00 263.76 12.66 ;
      LAYER Metal6 ;
        RECT 263.10 12.00 263.76 12.66 ;
      LAYER Metal3 ;
        RECT 263.10 12.00 263.76 12.66 ;
      LAYER Metal4 ;
        RECT 263.10 12.00 263.76 12.66 ;
    END
  END D1[19]
  PIN D1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 36.00 12.00 36.66 12.66 ;
      LAYER Metal6 ;
        RECT 36.00 12.00 36.66 12.66 ;
      LAYER Metal3 ;
        RECT 36.00 12.00 36.66 12.66 ;
      LAYER Metal4 ;
        RECT 36.00 12.00 36.66 12.66 ;
    END
  END D1[1]
  PIN D1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 264.24 12.00 264.90 12.66 ;
      LAYER Metal6 ;
        RECT 264.24 12.00 264.90 12.66 ;
      LAYER Metal3 ;
        RECT 264.24 12.00 264.90 12.66 ;
      LAYER Metal4 ;
        RECT 264.24 12.00 264.90 12.66 ;
    END
  END D1[20]
  PIN D1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 284.38 12.00 285.04 12.66 ;
      LAYER Metal6 ;
        RECT 284.38 12.00 285.04 12.66 ;
      LAYER Metal3 ;
        RECT 284.38 12.00 285.04 12.66 ;
      LAYER Metal4 ;
        RECT 284.38 12.00 285.04 12.66 ;
    END
  END D1[21]
  PIN D1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 285.52 12.00 286.18 12.66 ;
      LAYER Metal6 ;
        RECT 285.52 12.00 286.18 12.66 ;
      LAYER Metal3 ;
        RECT 285.52 12.00 286.18 12.66 ;
      LAYER Metal4 ;
        RECT 285.52 12.00 286.18 12.66 ;
    END
  END D1[22]
  PIN D1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 305.66 12.00 306.32 12.66 ;
      LAYER Metal6 ;
        RECT 305.66 12.00 306.32 12.66 ;
      LAYER Metal3 ;
        RECT 305.66 12.00 306.32 12.66 ;
      LAYER Metal4 ;
        RECT 305.66 12.00 306.32 12.66 ;
    END
  END D1[23]
  PIN D1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 306.80 12.00 307.46 12.66 ;
      LAYER Metal6 ;
        RECT 306.80 12.00 307.46 12.66 ;
      LAYER Metal3 ;
        RECT 306.80 12.00 307.46 12.66 ;
      LAYER Metal4 ;
        RECT 306.80 12.00 307.46 12.66 ;
    END
  END D1[24]
  PIN D1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 326.94 12.00 327.60 12.66 ;
      LAYER Metal6 ;
        RECT 326.94 12.00 327.60 12.66 ;
      LAYER Metal3 ;
        RECT 326.94 12.00 327.60 12.66 ;
      LAYER Metal4 ;
        RECT 326.94 12.00 327.60 12.66 ;
    END
  END D1[25]
  PIN D1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 328.08 12.00 328.74 12.66 ;
      LAYER Metal6 ;
        RECT 328.08 12.00 328.74 12.66 ;
      LAYER Metal3 ;
        RECT 328.08 12.00 328.74 12.66 ;
      LAYER Metal4 ;
        RECT 328.08 12.00 328.74 12.66 ;
    END
  END D1[26]
  PIN D1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 348.22 12.00 348.88 12.66 ;
      LAYER Metal6 ;
        RECT 348.22 12.00 348.88 12.66 ;
      LAYER Metal3 ;
        RECT 348.22 12.00 348.88 12.66 ;
      LAYER Metal4 ;
        RECT 348.22 12.00 348.88 12.66 ;
    END
  END D1[27]
  PIN D1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 349.36 12.00 350.02 12.66 ;
      LAYER Metal6 ;
        RECT 349.36 12.00 350.02 12.66 ;
      LAYER Metal3 ;
        RECT 349.36 12.00 350.02 12.66 ;
      LAYER Metal4 ;
        RECT 349.36 12.00 350.02 12.66 ;
    END
  END D1[28]
  PIN D1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 369.50 12.00 370.16 12.66 ;
      LAYER Metal6 ;
        RECT 369.50 12.00 370.16 12.66 ;
      LAYER Metal3 ;
        RECT 369.50 12.00 370.16 12.66 ;
      LAYER Metal4 ;
        RECT 369.50 12.00 370.16 12.66 ;
    END
  END D1[29]
  PIN D1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 37.14 12.00 37.80 12.66 ;
      LAYER Metal6 ;
        RECT 37.14 12.00 37.80 12.66 ;
      LAYER Metal3 ;
        RECT 37.14 12.00 37.80 12.66 ;
      LAYER Metal4 ;
        RECT 37.14 12.00 37.80 12.66 ;
    END
  END D1[2]
  PIN D1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 370.64 12.00 371.30 12.66 ;
      LAYER Metal6 ;
        RECT 370.64 12.00 371.30 12.66 ;
      LAYER Metal3 ;
        RECT 370.64 12.00 371.30 12.66 ;
      LAYER Metal4 ;
        RECT 370.64 12.00 371.30 12.66 ;
    END
  END D1[30]
  PIN D1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 390.78 12.00 391.44 12.66 ;
      LAYER Metal6 ;
        RECT 390.78 12.00 391.44 12.66 ;
      LAYER Metal3 ;
        RECT 390.78 12.00 391.44 12.66 ;
      LAYER Metal4 ;
        RECT 390.78 12.00 391.44 12.66 ;
    END
  END D1[31]
  PIN D1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 57.28 12.00 57.94 12.66 ;
      LAYER Metal6 ;
        RECT 57.28 12.00 57.94 12.66 ;
      LAYER Metal3 ;
        RECT 57.28 12.00 57.94 12.66 ;
      LAYER Metal4 ;
        RECT 57.28 12.00 57.94 12.66 ;
    END
  END D1[3]
  PIN D1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 58.42 12.00 59.08 12.66 ;
      LAYER Metal6 ;
        RECT 58.42 12.00 59.08 12.66 ;
      LAYER Metal3 ;
        RECT 58.42 12.00 59.08 12.66 ;
      LAYER Metal4 ;
        RECT 58.42 12.00 59.08 12.66 ;
    END
  END D1[4]
  PIN D1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 78.56 12.00 79.22 12.66 ;
      LAYER Metal6 ;
        RECT 78.56 12.00 79.22 12.66 ;
      LAYER Metal3 ;
        RECT 78.56 12.00 79.22 12.66 ;
      LAYER Metal4 ;
        RECT 78.56 12.00 79.22 12.66 ;
    END
  END D1[5]
  PIN D1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 79.70 12.00 80.36 12.66 ;
      LAYER Metal6 ;
        RECT 79.70 12.00 80.36 12.66 ;
      LAYER Metal3 ;
        RECT 79.70 12.00 80.36 12.66 ;
      LAYER Metal4 ;
        RECT 79.70 12.00 80.36 12.66 ;
    END
  END D1[6]
  PIN D1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 99.84 12.00 100.50 12.66 ;
      LAYER Metal6 ;
        RECT 99.84 12.00 100.50 12.66 ;
      LAYER Metal3 ;
        RECT 99.84 12.00 100.50 12.66 ;
      LAYER Metal4 ;
        RECT 99.84 12.00 100.50 12.66 ;
    END
  END D1[7]
  PIN D1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 100.98 12.00 101.64 12.66 ;
      LAYER Metal6 ;
        RECT 100.98 12.00 101.64 12.66 ;
      LAYER Metal3 ;
        RECT 100.98 12.00 101.64 12.66 ;
      LAYER Metal4 ;
        RECT 100.98 12.00 101.64 12.66 ;
    END
  END D1[8]
  PIN D1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 121.12 12.00 121.78 12.66 ;
      LAYER Metal6 ;
        RECT 121.12 12.00 121.78 12.66 ;
      LAYER Metal3 ;
        RECT 121.12 12.00 121.78 12.66 ;
      LAYER Metal4 ;
        RECT 121.12 12.00 121.78 12.66 ;
    END
  END D1[9]
  PIN D2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 25.36 12.00 26.02 12.66 ;
      LAYER Metal6 ;
        RECT 25.36 12.00 26.02 12.66 ;
      LAYER Metal3 ;
        RECT 25.36 12.00 26.02 12.66 ;
      LAYER Metal4 ;
        RECT 25.36 12.00 26.02 12.66 ;
    END
  END D2[0]
  PIN D2[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 131.76 12.00 132.42 12.66 ;
      LAYER Metal6 ;
        RECT 131.76 12.00 132.42 12.66 ;
      LAYER Metal3 ;
        RECT 131.76 12.00 132.42 12.66 ;
      LAYER Metal4 ;
        RECT 131.76 12.00 132.42 12.66 ;
    END
  END D2[10]
  PIN D2[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 132.90 12.00 133.56 12.66 ;
      LAYER Metal6 ;
        RECT 132.90 12.00 133.56 12.66 ;
      LAYER Metal3 ;
        RECT 132.90 12.00 133.56 12.66 ;
      LAYER Metal4 ;
        RECT 132.90 12.00 133.56 12.66 ;
    END
  END D2[11]
  PIN D2[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 153.04 12.00 153.70 12.66 ;
      LAYER Metal6 ;
        RECT 153.04 12.00 153.70 12.66 ;
      LAYER Metal3 ;
        RECT 153.04 12.00 153.70 12.66 ;
      LAYER Metal4 ;
        RECT 153.04 12.00 153.70 12.66 ;
    END
  END D2[12]
  PIN D2[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 154.18 12.00 154.84 12.66 ;
      LAYER Metal6 ;
        RECT 154.18 12.00 154.84 12.66 ;
      LAYER Metal3 ;
        RECT 154.18 12.00 154.84 12.66 ;
      LAYER Metal4 ;
        RECT 154.18 12.00 154.84 12.66 ;
    END
  END D2[13]
  PIN D2[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 174.32 12.00 174.98 12.66 ;
      LAYER Metal6 ;
        RECT 174.32 12.00 174.98 12.66 ;
      LAYER Metal3 ;
        RECT 174.32 12.00 174.98 12.66 ;
      LAYER Metal4 ;
        RECT 174.32 12.00 174.98 12.66 ;
    END
  END D2[14]
  PIN D2[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 175.46 12.00 176.12 12.66 ;
      LAYER Metal6 ;
        RECT 175.46 12.00 176.12 12.66 ;
      LAYER Metal3 ;
        RECT 175.46 12.00 176.12 12.66 ;
      LAYER Metal4 ;
        RECT 175.46 12.00 176.12 12.66 ;
    END
  END D2[15]
  PIN D2[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 231.18 12.00 231.84 12.66 ;
      LAYER Metal6 ;
        RECT 231.18 12.00 231.84 12.66 ;
      LAYER Metal3 ;
        RECT 231.18 12.00 231.84 12.66 ;
      LAYER Metal4 ;
        RECT 231.18 12.00 231.84 12.66 ;
    END
  END D2[16]
  PIN D2[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 232.32 12.00 232.98 12.66 ;
      LAYER Metal6 ;
        RECT 232.32 12.00 232.98 12.66 ;
      LAYER Metal3 ;
        RECT 232.32 12.00 232.98 12.66 ;
      LAYER Metal4 ;
        RECT 232.32 12.00 232.98 12.66 ;
    END
  END D2[17]
  PIN D2[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 252.46 12.00 253.12 12.66 ;
      LAYER Metal6 ;
        RECT 252.46 12.00 253.12 12.66 ;
      LAYER Metal3 ;
        RECT 252.46 12.00 253.12 12.66 ;
      LAYER Metal4 ;
        RECT 252.46 12.00 253.12 12.66 ;
    END
  END D2[18]
  PIN D2[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 253.60 12.00 254.26 12.66 ;
      LAYER Metal6 ;
        RECT 253.60 12.00 254.26 12.66 ;
      LAYER Metal3 ;
        RECT 253.60 12.00 254.26 12.66 ;
      LAYER Metal4 ;
        RECT 253.60 12.00 254.26 12.66 ;
    END
  END D2[19]
  PIN D2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 26.50 12.00 27.16 12.66 ;
      LAYER Metal6 ;
        RECT 26.50 12.00 27.16 12.66 ;
      LAYER Metal3 ;
        RECT 26.50 12.00 27.16 12.66 ;
      LAYER Metal4 ;
        RECT 26.50 12.00 27.16 12.66 ;
    END
  END D2[1]
  PIN D2[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 273.74 12.00 274.40 12.66 ;
      LAYER Metal6 ;
        RECT 273.74 12.00 274.40 12.66 ;
      LAYER Metal3 ;
        RECT 273.74 12.00 274.40 12.66 ;
      LAYER Metal4 ;
        RECT 273.74 12.00 274.40 12.66 ;
    END
  END D2[20]
  PIN D2[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 274.88 12.00 275.54 12.66 ;
      LAYER Metal6 ;
        RECT 274.88 12.00 275.54 12.66 ;
      LAYER Metal3 ;
        RECT 274.88 12.00 275.54 12.66 ;
      LAYER Metal4 ;
        RECT 274.88 12.00 275.54 12.66 ;
    END
  END D2[21]
  PIN D2[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 295.02 12.00 295.68 12.66 ;
      LAYER Metal6 ;
        RECT 295.02 12.00 295.68 12.66 ;
      LAYER Metal3 ;
        RECT 295.02 12.00 295.68 12.66 ;
      LAYER Metal4 ;
        RECT 295.02 12.00 295.68 12.66 ;
    END
  END D2[22]
  PIN D2[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 296.16 12.00 296.82 12.66 ;
      LAYER Metal6 ;
        RECT 296.16 12.00 296.82 12.66 ;
      LAYER Metal3 ;
        RECT 296.16 12.00 296.82 12.66 ;
      LAYER Metal4 ;
        RECT 296.16 12.00 296.82 12.66 ;
    END
  END D2[23]
  PIN D2[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 316.30 12.00 316.96 12.66 ;
      LAYER Metal6 ;
        RECT 316.30 12.00 316.96 12.66 ;
      LAYER Metal3 ;
        RECT 316.30 12.00 316.96 12.66 ;
      LAYER Metal4 ;
        RECT 316.30 12.00 316.96 12.66 ;
    END
  END D2[24]
  PIN D2[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 317.44 12.00 318.10 12.66 ;
      LAYER Metal6 ;
        RECT 317.44 12.00 318.10 12.66 ;
      LAYER Metal3 ;
        RECT 317.44 12.00 318.10 12.66 ;
      LAYER Metal4 ;
        RECT 317.44 12.00 318.10 12.66 ;
    END
  END D2[25]
  PIN D2[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 337.58 12.00 338.24 12.66 ;
      LAYER Metal6 ;
        RECT 337.58 12.00 338.24 12.66 ;
      LAYER Metal3 ;
        RECT 337.58 12.00 338.24 12.66 ;
      LAYER Metal4 ;
        RECT 337.58 12.00 338.24 12.66 ;
    END
  END D2[26]
  PIN D2[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 338.72 12.00 339.38 12.66 ;
      LAYER Metal6 ;
        RECT 338.72 12.00 339.38 12.66 ;
      LAYER Metal3 ;
        RECT 338.72 12.00 339.38 12.66 ;
      LAYER Metal4 ;
        RECT 338.72 12.00 339.38 12.66 ;
    END
  END D2[27]
  PIN D2[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 358.86 12.00 359.52 12.66 ;
      LAYER Metal6 ;
        RECT 358.86 12.00 359.52 12.66 ;
      LAYER Metal3 ;
        RECT 358.86 12.00 359.52 12.66 ;
      LAYER Metal4 ;
        RECT 358.86 12.00 359.52 12.66 ;
    END
  END D2[28]
  PIN D2[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 360.00 12.00 360.66 12.66 ;
      LAYER Metal6 ;
        RECT 360.00 12.00 360.66 12.66 ;
      LAYER Metal3 ;
        RECT 360.00 12.00 360.66 12.66 ;
      LAYER Metal4 ;
        RECT 360.00 12.00 360.66 12.66 ;
    END
  END D2[29]
  PIN D2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 46.64 12.00 47.30 12.66 ;
      LAYER Metal6 ;
        RECT 46.64 12.00 47.30 12.66 ;
      LAYER Metal3 ;
        RECT 46.64 12.00 47.30 12.66 ;
      LAYER Metal4 ;
        RECT 46.64 12.00 47.30 12.66 ;
    END
  END D2[2]
  PIN D2[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 380.14 12.00 380.80 12.66 ;
      LAYER Metal6 ;
        RECT 380.14 12.00 380.80 12.66 ;
      LAYER Metal3 ;
        RECT 380.14 12.00 380.80 12.66 ;
      LAYER Metal4 ;
        RECT 380.14 12.00 380.80 12.66 ;
    END
  END D2[30]
  PIN D2[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 381.28 12.00 381.94 12.66 ;
      LAYER Metal6 ;
        RECT 381.28 12.00 381.94 12.66 ;
      LAYER Metal3 ;
        RECT 381.28 12.00 381.94 12.66 ;
      LAYER Metal4 ;
        RECT 381.28 12.00 381.94 12.66 ;
    END
  END D2[31]
  PIN D2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 47.78 12.00 48.44 12.66 ;
      LAYER Metal6 ;
        RECT 47.78 12.00 48.44 12.66 ;
      LAYER Metal3 ;
        RECT 47.78 12.00 48.44 12.66 ;
      LAYER Metal4 ;
        RECT 47.78 12.00 48.44 12.66 ;
    END
  END D2[3]
  PIN D2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 67.92 12.00 68.58 12.66 ;
      LAYER Metal6 ;
        RECT 67.92 12.00 68.58 12.66 ;
      LAYER Metal3 ;
        RECT 67.92 12.00 68.58 12.66 ;
      LAYER Metal4 ;
        RECT 67.92 12.00 68.58 12.66 ;
    END
  END D2[4]
  PIN D2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 69.06 12.00 69.72 12.66 ;
      LAYER Metal6 ;
        RECT 69.06 12.00 69.72 12.66 ;
      LAYER Metal3 ;
        RECT 69.06 12.00 69.72 12.66 ;
      LAYER Metal4 ;
        RECT 69.06 12.00 69.72 12.66 ;
    END
  END D2[5]
  PIN D2[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 89.20 12.00 89.86 12.66 ;
      LAYER Metal6 ;
        RECT 89.20 12.00 89.86 12.66 ;
      LAYER Metal3 ;
        RECT 89.20 12.00 89.86 12.66 ;
      LAYER Metal4 ;
        RECT 89.20 12.00 89.86 12.66 ;
    END
  END D2[6]
  PIN D2[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 90.34 12.00 91.00 12.66 ;
      LAYER Metal6 ;
        RECT 90.34 12.00 91.00 12.66 ;
      LAYER Metal3 ;
        RECT 90.34 12.00 91.00 12.66 ;
      LAYER Metal4 ;
        RECT 90.34 12.00 91.00 12.66 ;
    END
  END D2[7]
  PIN D2[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 110.48 12.00 111.14 12.66 ;
      LAYER Metal6 ;
        RECT 110.48 12.00 111.14 12.66 ;
      LAYER Metal3 ;
        RECT 110.48 12.00 111.14 12.66 ;
      LAYER Metal4 ;
        RECT 110.48 12.00 111.14 12.66 ;
    END
  END D2[8]
  PIN D2[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 111.62 12.00 112.28 12.66 ;
      LAYER Metal6 ;
        RECT 111.62 12.00 112.28 12.66 ;
      LAYER Metal3 ;
        RECT 111.62 12.00 112.28 12.66 ;
      LAYER Metal4 ;
        RECT 111.62 12.00 112.28 12.66 ;
    END
  END D2[9]
  PIN Q1[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 18.28 12.00 18.94 12.66 ;
      LAYER Metal6 ;
        RECT 18.28 12.00 18.94 12.66 ;
      LAYER Metal3 ;
        RECT 18.28 12.00 18.94 12.66 ;
      LAYER Metal4 ;
        RECT 18.28 12.00 18.94 12.66 ;
    END
  END Q1[0]
  PIN Q1[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 125.56 12.00 126.22 12.66 ;
      LAYER Metal6 ;
        RECT 125.56 12.00 126.22 12.66 ;
      LAYER Metal3 ;
        RECT 125.56 12.00 126.22 12.66 ;
      LAYER Metal4 ;
        RECT 125.56 12.00 126.22 12.66 ;
    END
  END Q1[10]
  PIN Q1[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 139.10 12.00 139.76 12.66 ;
      LAYER Metal6 ;
        RECT 139.10 12.00 139.76 12.66 ;
      LAYER Metal3 ;
        RECT 139.10 12.00 139.76 12.66 ;
      LAYER Metal4 ;
        RECT 139.10 12.00 139.76 12.66 ;
    END
  END Q1[11]
  PIN Q1[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 146.84 12.00 147.50 12.66 ;
      LAYER Metal6 ;
        RECT 146.84 12.00 147.50 12.66 ;
      LAYER Metal3 ;
        RECT 146.84 12.00 147.50 12.66 ;
      LAYER Metal4 ;
        RECT 146.84 12.00 147.50 12.66 ;
    END
  END Q1[12]
  PIN Q1[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 160.38 12.00 161.04 12.66 ;
      LAYER Metal6 ;
        RECT 160.38 12.00 161.04 12.66 ;
      LAYER Metal3 ;
        RECT 160.38 12.00 161.04 12.66 ;
      LAYER Metal4 ;
        RECT 160.38 12.00 161.04 12.66 ;
    END
  END Q1[13]
  PIN Q1[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 168.12 12.00 168.78 12.66 ;
      LAYER Metal6 ;
        RECT 168.12 12.00 168.78 12.66 ;
      LAYER Metal3 ;
        RECT 168.12 12.00 168.78 12.66 ;
      LAYER Metal4 ;
        RECT 168.12 12.00 168.78 12.66 ;
    END
  END Q1[14]
  PIN Q1[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 181.66 12.00 182.32 12.66 ;
      LAYER Metal6 ;
        RECT 181.66 12.00 182.32 12.66 ;
      LAYER Metal3 ;
        RECT 181.66 12.00 182.32 12.66 ;
      LAYER Metal4 ;
        RECT 181.66 12.00 182.32 12.66 ;
    END
  END Q1[15]
  PIN Q1[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 224.98 12.00 225.64 12.66 ;
      LAYER Metal6 ;
        RECT 224.98 12.00 225.64 12.66 ;
      LAYER Metal3 ;
        RECT 224.98 12.00 225.64 12.66 ;
      LAYER Metal4 ;
        RECT 224.98 12.00 225.64 12.66 ;
    END
  END Q1[16]
  PIN Q1[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 238.52 12.00 239.18 12.66 ;
      LAYER Metal6 ;
        RECT 238.52 12.00 239.18 12.66 ;
      LAYER Metal3 ;
        RECT 238.52 12.00 239.18 12.66 ;
      LAYER Metal4 ;
        RECT 238.52 12.00 239.18 12.66 ;
    END
  END Q1[17]
  PIN Q1[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 246.26 12.00 246.92 12.66 ;
      LAYER Metal6 ;
        RECT 246.26 12.00 246.92 12.66 ;
      LAYER Metal3 ;
        RECT 246.26 12.00 246.92 12.66 ;
      LAYER Metal4 ;
        RECT 246.26 12.00 246.92 12.66 ;
    END
  END Q1[18]
  PIN Q1[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 259.80 12.00 260.46 12.66 ;
      LAYER Metal6 ;
        RECT 259.80 12.00 260.46 12.66 ;
      LAYER Metal3 ;
        RECT 259.80 12.00 260.46 12.66 ;
      LAYER Metal4 ;
        RECT 259.80 12.00 260.46 12.66 ;
    END
  END Q1[19]
  PIN Q1[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 32.70 12.00 33.36 12.66 ;
      LAYER Metal6 ;
        RECT 32.70 12.00 33.36 12.66 ;
      LAYER Metal3 ;
        RECT 32.70 12.00 33.36 12.66 ;
      LAYER Metal4 ;
        RECT 32.70 12.00 33.36 12.66 ;
    END
  END Q1[1]
  PIN Q1[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 267.54 12.00 268.20 12.66 ;
      LAYER Metal6 ;
        RECT 267.54 12.00 268.20 12.66 ;
      LAYER Metal3 ;
        RECT 267.54 12.00 268.20 12.66 ;
      LAYER Metal4 ;
        RECT 267.54 12.00 268.20 12.66 ;
    END
  END Q1[20]
  PIN Q1[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 281.08 12.00 281.74 12.66 ;
      LAYER Metal6 ;
        RECT 281.08 12.00 281.74 12.66 ;
      LAYER Metal3 ;
        RECT 281.08 12.00 281.74 12.66 ;
      LAYER Metal4 ;
        RECT 281.08 12.00 281.74 12.66 ;
    END
  END Q1[21]
  PIN Q1[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 288.82 12.00 289.48 12.66 ;
      LAYER Metal6 ;
        RECT 288.82 12.00 289.48 12.66 ;
      LAYER Metal3 ;
        RECT 288.82 12.00 289.48 12.66 ;
      LAYER Metal4 ;
        RECT 288.82 12.00 289.48 12.66 ;
    END
  END Q1[22]
  PIN Q1[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 302.36 12.00 303.02 12.66 ;
      LAYER Metal6 ;
        RECT 302.36 12.00 303.02 12.66 ;
      LAYER Metal3 ;
        RECT 302.36 12.00 303.02 12.66 ;
      LAYER Metal4 ;
        RECT 302.36 12.00 303.02 12.66 ;
    END
  END Q1[23]
  PIN Q1[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 310.10 12.00 310.76 12.66 ;
      LAYER Metal6 ;
        RECT 310.10 12.00 310.76 12.66 ;
      LAYER Metal3 ;
        RECT 310.10 12.00 310.76 12.66 ;
      LAYER Metal4 ;
        RECT 310.10 12.00 310.76 12.66 ;
    END
  END Q1[24]
  PIN Q1[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 323.64 12.00 324.30 12.66 ;
      LAYER Metal6 ;
        RECT 323.64 12.00 324.30 12.66 ;
      LAYER Metal3 ;
        RECT 323.64 12.00 324.30 12.66 ;
      LAYER Metal4 ;
        RECT 323.64 12.00 324.30 12.66 ;
    END
  END Q1[25]
  PIN Q1[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 331.38 12.00 332.04 12.66 ;
      LAYER Metal6 ;
        RECT 331.38 12.00 332.04 12.66 ;
      LAYER Metal3 ;
        RECT 331.38 12.00 332.04 12.66 ;
      LAYER Metal4 ;
        RECT 331.38 12.00 332.04 12.66 ;
    END
  END Q1[26]
  PIN Q1[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 344.92 12.00 345.58 12.66 ;
      LAYER Metal6 ;
        RECT 344.92 12.00 345.58 12.66 ;
      LAYER Metal3 ;
        RECT 344.92 12.00 345.58 12.66 ;
      LAYER Metal4 ;
        RECT 344.92 12.00 345.58 12.66 ;
    END
  END Q1[27]
  PIN Q1[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 352.66 12.00 353.32 12.66 ;
      LAYER Metal6 ;
        RECT 352.66 12.00 353.32 12.66 ;
      LAYER Metal3 ;
        RECT 352.66 12.00 353.32 12.66 ;
      LAYER Metal4 ;
        RECT 352.66 12.00 353.32 12.66 ;
    END
  END Q1[28]
  PIN Q1[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 366.20 12.00 366.86 12.66 ;
      LAYER Metal6 ;
        RECT 366.20 12.00 366.86 12.66 ;
      LAYER Metal3 ;
        RECT 366.20 12.00 366.86 12.66 ;
      LAYER Metal4 ;
        RECT 366.20 12.00 366.86 12.66 ;
    END
  END Q1[29]
  PIN Q1[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 40.44 12.00 41.10 12.66 ;
      LAYER Metal6 ;
        RECT 40.44 12.00 41.10 12.66 ;
      LAYER Metal3 ;
        RECT 40.44 12.00 41.10 12.66 ;
      LAYER Metal4 ;
        RECT 40.44 12.00 41.10 12.66 ;
    END
  END Q1[2]
  PIN Q1[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 373.94 12.00 374.60 12.66 ;
      LAYER Metal6 ;
        RECT 373.94 12.00 374.60 12.66 ;
      LAYER Metal3 ;
        RECT 373.94 12.00 374.60 12.66 ;
      LAYER Metal4 ;
        RECT 373.94 12.00 374.60 12.66 ;
    END
  END Q1[30]
  PIN Q1[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 388.36 12.00 389.02 12.66 ;
      LAYER Metal6 ;
        RECT 388.36 12.00 389.02 12.66 ;
      LAYER Metal3 ;
        RECT 388.36 12.00 389.02 12.66 ;
      LAYER Metal4 ;
        RECT 388.36 12.00 389.02 12.66 ;
    END
  END Q1[31]
  PIN Q1[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 53.98 12.00 54.64 12.66 ;
      LAYER Metal6 ;
        RECT 53.98 12.00 54.64 12.66 ;
      LAYER Metal3 ;
        RECT 53.98 12.00 54.64 12.66 ;
      LAYER Metal4 ;
        RECT 53.98 12.00 54.64 12.66 ;
    END
  END Q1[3]
  PIN Q1[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 61.72 12.00 62.38 12.66 ;
      LAYER Metal6 ;
        RECT 61.72 12.00 62.38 12.66 ;
      LAYER Metal3 ;
        RECT 61.72 12.00 62.38 12.66 ;
      LAYER Metal4 ;
        RECT 61.72 12.00 62.38 12.66 ;
    END
  END Q1[4]
  PIN Q1[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 75.26 12.00 75.92 12.66 ;
      LAYER Metal6 ;
        RECT 75.26 12.00 75.92 12.66 ;
      LAYER Metal3 ;
        RECT 75.26 12.00 75.92 12.66 ;
      LAYER Metal4 ;
        RECT 75.26 12.00 75.92 12.66 ;
    END
  END Q1[5]
  PIN Q1[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 83.00 12.00 83.66 12.66 ;
      LAYER Metal6 ;
        RECT 83.00 12.00 83.66 12.66 ;
      LAYER Metal3 ;
        RECT 83.00 12.00 83.66 12.66 ;
      LAYER Metal4 ;
        RECT 83.00 12.00 83.66 12.66 ;
    END
  END Q1[6]
  PIN Q1[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 96.54 12.00 97.20 12.66 ;
      LAYER Metal6 ;
        RECT 96.54 12.00 97.20 12.66 ;
      LAYER Metal3 ;
        RECT 96.54 12.00 97.20 12.66 ;
      LAYER Metal4 ;
        RECT 96.54 12.00 97.20 12.66 ;
    END
  END Q1[7]
  PIN Q1[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 104.28 12.00 104.94 12.66 ;
      LAYER Metal6 ;
        RECT 104.28 12.00 104.94 12.66 ;
      LAYER Metal3 ;
        RECT 104.28 12.00 104.94 12.66 ;
      LAYER Metal4 ;
        RECT 104.28 12.00 104.94 12.66 ;
    END
  END Q1[8]
  PIN Q1[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 117.82 12.00 118.48 12.66 ;
      LAYER Metal6 ;
        RECT 117.82 12.00 118.48 12.66 ;
      LAYER Metal3 ;
        RECT 117.82 12.00 118.48 12.66 ;
      LAYER Metal4 ;
        RECT 117.82 12.00 118.48 12.66 ;
    END
  END Q1[9]
  PIN Q2[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 22.06 12.00 22.72 12.66 ;
      LAYER Metal6 ;
        RECT 22.06 12.00 22.72 12.66 ;
      LAYER Metal3 ;
        RECT 22.06 12.00 22.72 12.66 ;
      LAYER Metal4 ;
        RECT 22.06 12.00 22.72 12.66 ;
    END
  END Q2[0]
  PIN Q2[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 128.46 12.00 129.12 12.66 ;
      LAYER Metal6 ;
        RECT 128.46 12.00 129.12 12.66 ;
      LAYER Metal3 ;
        RECT 128.46 12.00 129.12 12.66 ;
      LAYER Metal4 ;
        RECT 128.46 12.00 129.12 12.66 ;
    END
  END Q2[10]
  PIN Q2[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 136.20 12.00 136.86 12.66 ;
      LAYER Metal6 ;
        RECT 136.20 12.00 136.86 12.66 ;
      LAYER Metal3 ;
        RECT 136.20 12.00 136.86 12.66 ;
      LAYER Metal4 ;
        RECT 136.20 12.00 136.86 12.66 ;
    END
  END Q2[11]
  PIN Q2[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 149.74 12.00 150.40 12.66 ;
      LAYER Metal6 ;
        RECT 149.74 12.00 150.40 12.66 ;
      LAYER Metal3 ;
        RECT 149.74 12.00 150.40 12.66 ;
      LAYER Metal4 ;
        RECT 149.74 12.00 150.40 12.66 ;
    END
  END Q2[12]
  PIN Q2[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 157.48 12.00 158.14 12.66 ;
      LAYER Metal6 ;
        RECT 157.48 12.00 158.14 12.66 ;
      LAYER Metal3 ;
        RECT 157.48 12.00 158.14 12.66 ;
      LAYER Metal4 ;
        RECT 157.48 12.00 158.14 12.66 ;
    END
  END Q2[13]
  PIN Q2[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 171.02 12.00 171.68 12.66 ;
      LAYER Metal6 ;
        RECT 171.02 12.00 171.68 12.66 ;
      LAYER Metal3 ;
        RECT 171.02 12.00 171.68 12.66 ;
      LAYER Metal4 ;
        RECT 171.02 12.00 171.68 12.66 ;
    END
  END Q2[14]
  PIN Q2[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 178.76 12.00 179.42 12.66 ;
      LAYER Metal6 ;
        RECT 178.76 12.00 179.42 12.66 ;
      LAYER Metal3 ;
        RECT 178.76 12.00 179.42 12.66 ;
      LAYER Metal4 ;
        RECT 178.76 12.00 179.42 12.66 ;
    END
  END Q2[15]
  PIN Q2[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 227.88 12.00 228.54 12.66 ;
      LAYER Metal6 ;
        RECT 227.88 12.00 228.54 12.66 ;
      LAYER Metal3 ;
        RECT 227.88 12.00 228.54 12.66 ;
      LAYER Metal4 ;
        RECT 227.88 12.00 228.54 12.66 ;
    END
  END Q2[16]
  PIN Q2[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 235.62 12.00 236.28 12.66 ;
      LAYER Metal6 ;
        RECT 235.62 12.00 236.28 12.66 ;
      LAYER Metal3 ;
        RECT 235.62 12.00 236.28 12.66 ;
      LAYER Metal4 ;
        RECT 235.62 12.00 236.28 12.66 ;
    END
  END Q2[17]
  PIN Q2[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 249.16 12.00 249.82 12.66 ;
      LAYER Metal6 ;
        RECT 249.16 12.00 249.82 12.66 ;
      LAYER Metal3 ;
        RECT 249.16 12.00 249.82 12.66 ;
      LAYER Metal4 ;
        RECT 249.16 12.00 249.82 12.66 ;
    END
  END Q2[18]
  PIN Q2[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 256.90 12.00 257.56 12.66 ;
      LAYER Metal6 ;
        RECT 256.90 12.00 257.56 12.66 ;
      LAYER Metal3 ;
        RECT 256.90 12.00 257.56 12.66 ;
      LAYER Metal4 ;
        RECT 256.90 12.00 257.56 12.66 ;
    END
  END Q2[19]
  PIN Q2[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 29.80 12.00 30.46 12.66 ;
      LAYER Metal6 ;
        RECT 29.80 12.00 30.46 12.66 ;
      LAYER Metal3 ;
        RECT 29.80 12.00 30.46 12.66 ;
      LAYER Metal4 ;
        RECT 29.80 12.00 30.46 12.66 ;
    END
  END Q2[1]
  PIN Q2[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 270.44 12.00 271.10 12.66 ;
      LAYER Metal6 ;
        RECT 270.44 12.00 271.10 12.66 ;
      LAYER Metal3 ;
        RECT 270.44 12.00 271.10 12.66 ;
      LAYER Metal4 ;
        RECT 270.44 12.00 271.10 12.66 ;
    END
  END Q2[20]
  PIN Q2[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 278.18 12.00 278.84 12.66 ;
      LAYER Metal6 ;
        RECT 278.18 12.00 278.84 12.66 ;
      LAYER Metal3 ;
        RECT 278.18 12.00 278.84 12.66 ;
      LAYER Metal4 ;
        RECT 278.18 12.00 278.84 12.66 ;
    END
  END Q2[21]
  PIN Q2[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 291.72 12.00 292.38 12.66 ;
      LAYER Metal6 ;
        RECT 291.72 12.00 292.38 12.66 ;
      LAYER Metal3 ;
        RECT 291.72 12.00 292.38 12.66 ;
      LAYER Metal4 ;
        RECT 291.72 12.00 292.38 12.66 ;
    END
  END Q2[22]
  PIN Q2[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 299.46 12.00 300.12 12.66 ;
      LAYER Metal6 ;
        RECT 299.46 12.00 300.12 12.66 ;
      LAYER Metal3 ;
        RECT 299.46 12.00 300.12 12.66 ;
      LAYER Metal4 ;
        RECT 299.46 12.00 300.12 12.66 ;
    END
  END Q2[23]
  PIN Q2[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 313.00 12.00 313.66 12.66 ;
      LAYER Metal6 ;
        RECT 313.00 12.00 313.66 12.66 ;
      LAYER Metal3 ;
        RECT 313.00 12.00 313.66 12.66 ;
      LAYER Metal4 ;
        RECT 313.00 12.00 313.66 12.66 ;
    END
  END Q2[24]
  PIN Q2[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 320.74 12.00 321.40 12.66 ;
      LAYER Metal6 ;
        RECT 320.74 12.00 321.40 12.66 ;
      LAYER Metal3 ;
        RECT 320.74 12.00 321.40 12.66 ;
      LAYER Metal4 ;
        RECT 320.74 12.00 321.40 12.66 ;
    END
  END Q2[25]
  PIN Q2[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 334.28 12.00 334.94 12.66 ;
      LAYER Metal6 ;
        RECT 334.28 12.00 334.94 12.66 ;
      LAYER Metal3 ;
        RECT 334.28 12.00 334.94 12.66 ;
      LAYER Metal4 ;
        RECT 334.28 12.00 334.94 12.66 ;
    END
  END Q2[26]
  PIN Q2[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 342.02 12.00 342.68 12.66 ;
      LAYER Metal6 ;
        RECT 342.02 12.00 342.68 12.66 ;
      LAYER Metal3 ;
        RECT 342.02 12.00 342.68 12.66 ;
      LAYER Metal4 ;
        RECT 342.02 12.00 342.68 12.66 ;
    END
  END Q2[27]
  PIN Q2[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 355.56 12.00 356.22 12.66 ;
      LAYER Metal6 ;
        RECT 355.56 12.00 356.22 12.66 ;
      LAYER Metal3 ;
        RECT 355.56 12.00 356.22 12.66 ;
      LAYER Metal4 ;
        RECT 355.56 12.00 356.22 12.66 ;
    END
  END Q2[28]
  PIN Q2[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 363.30 12.00 363.96 12.66 ;
      LAYER Metal6 ;
        RECT 363.30 12.00 363.96 12.66 ;
      LAYER Metal3 ;
        RECT 363.30 12.00 363.96 12.66 ;
      LAYER Metal4 ;
        RECT 363.30 12.00 363.96 12.66 ;
    END
  END Q2[29]
  PIN Q2[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 43.34 12.00 44.00 12.66 ;
      LAYER Metal6 ;
        RECT 43.34 12.00 44.00 12.66 ;
      LAYER Metal3 ;
        RECT 43.34 12.00 44.00 12.66 ;
      LAYER Metal4 ;
        RECT 43.34 12.00 44.00 12.66 ;
    END
  END Q2[2]
  PIN Q2[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 376.84 12.00 377.50 12.66 ;
      LAYER Metal6 ;
        RECT 376.84 12.00 377.50 12.66 ;
      LAYER Metal3 ;
        RECT 376.84 12.00 377.50 12.66 ;
      LAYER Metal4 ;
        RECT 376.84 12.00 377.50 12.66 ;
    END
  END Q2[30]
  PIN Q2[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 384.58 12.00 385.24 12.66 ;
      LAYER Metal6 ;
        RECT 384.58 12.00 385.24 12.66 ;
      LAYER Metal3 ;
        RECT 384.58 12.00 385.24 12.66 ;
      LAYER Metal4 ;
        RECT 384.58 12.00 385.24 12.66 ;
    END
  END Q2[31]
  PIN Q2[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 51.08 12.00 51.74 12.66 ;
      LAYER Metal6 ;
        RECT 51.08 12.00 51.74 12.66 ;
      LAYER Metal3 ;
        RECT 51.08 12.00 51.74 12.66 ;
      LAYER Metal4 ;
        RECT 51.08 12.00 51.74 12.66 ;
    END
  END Q2[3]
  PIN Q2[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 64.62 12.00 65.28 12.66 ;
      LAYER Metal6 ;
        RECT 64.62 12.00 65.28 12.66 ;
      LAYER Metal3 ;
        RECT 64.62 12.00 65.28 12.66 ;
      LAYER Metal4 ;
        RECT 64.62 12.00 65.28 12.66 ;
    END
  END Q2[4]
  PIN Q2[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 72.36 12.00 73.02 12.66 ;
      LAYER Metal6 ;
        RECT 72.36 12.00 73.02 12.66 ;
      LAYER Metal3 ;
        RECT 72.36 12.00 73.02 12.66 ;
      LAYER Metal4 ;
        RECT 72.36 12.00 73.02 12.66 ;
    END
  END Q2[5]
  PIN Q2[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 85.90 12.00 86.56 12.66 ;
      LAYER Metal6 ;
        RECT 85.90 12.00 86.56 12.66 ;
      LAYER Metal3 ;
        RECT 85.90 12.00 86.56 12.66 ;
      LAYER Metal4 ;
        RECT 85.90 12.00 86.56 12.66 ;
    END
  END Q2[6]
  PIN Q2[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 93.64 12.00 94.30 12.66 ;
      LAYER Metal6 ;
        RECT 93.64 12.00 94.30 12.66 ;
      LAYER Metal3 ;
        RECT 93.64 12.00 94.30 12.66 ;
      LAYER Metal4 ;
        RECT 93.64 12.00 94.30 12.66 ;
    END
  END Q2[7]
  PIN Q2[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 107.18 12.00 107.84 12.66 ;
      LAYER Metal6 ;
        RECT 107.18 12.00 107.84 12.66 ;
      LAYER Metal3 ;
        RECT 107.18 12.00 107.84 12.66 ;
      LAYER Metal4 ;
        RECT 107.18 12.00 107.84 12.66 ;
    END
  END Q2[8]
  PIN Q2[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 114.92 12.00 115.58 12.66 ;
      LAYER Metal6 ;
        RECT 114.92 12.00 115.58 12.66 ;
      LAYER Metal3 ;
        RECT 114.92 12.00 115.58 12.66 ;
      LAYER Metal4 ;
        RECT 114.92 12.00 115.58 12.66 ;
    END
  END Q2[9]
  PIN WE1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 212.68 12.00 213.34 12.66 ;
      LAYER Metal6 ;
        RECT 212.68 12.00 213.34 12.66 ;
      LAYER Metal3 ;
        RECT 212.68 12.00 213.34 12.66 ;
      LAYER Metal4 ;
        RECT 212.68 12.00 213.34 12.66 ;
    END
  END WE1
  PIN WE2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 193.96 12.00 194.62 12.66 ;
      LAYER Metal6 ;
        RECT 193.96 12.00 194.62 12.66 ;
      LAYER Metal3 ;
        RECT 193.96 12.00 194.62 12.66 ;
      LAYER Metal4 ;
        RECT 193.96 12.00 194.62 12.66 ;
    END
  END WE2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE RING ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 140.03 423.01 145.03 ;
        RECT 0.00 0.00 423.01 5.00 ;
      LAYER Metal2 ;
        RECT 418.01 0.00 423.01 145.03 ;
        RECT 0.00 0.00 5.00 145.03 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE RING ;
    PORT
      LAYER Metal1 ;
        RECT 5.60 134.44 417.42 139.44 ;
        RECT 5.60 5.60 417.42 10.60 ;
      LAYER Metal2 ;
        RECT 412.42 5.60 417.42 139.44 ;
        RECT 5.60 5.60 10.60 139.44 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      RECT 12.00 12.00 411.02 132.97 ;
    LAYER Metal2 ;
      RECT 12.00 12.00 411.02 132.97 ;
    LAYER Metal3 ;
#      RECT 12.00 12.00 411.02 132.97 ;
        RECT 12.84 12.84 411.02 132.97 ;
        RECT 12.00 12.00 15.68 36.22 ;
        RECT 16.70 12.00 18.10 132.97 ;
        RECT 19.12 12.00 21.88 132.97 ;
        RECT 22.90 12.00 25.18 132.97 ;
        RECT 26.20 12.00 26.32 132.97 ;
        RECT 27.34 12.00 29.62 132.97 ;
        RECT 30.64 12.00 32.52 132.97 ;
        RECT 33.54 12.00 35.82 132.97 ;
        RECT 36.84 12.00 36.96 132.97 ;
        RECT 37.98 12.00 40.26 132.97 ;
        RECT 41.28 12.00 43.16 132.97 ;
        RECT 44.18 12.00 46.46 132.97 ;
        RECT 47.48 12.00 47.60 132.97 ;
        RECT 48.62 12.00 50.90 132.97 ;
        RECT 51.92 12.00 53.80 132.97 ;
        RECT 54.82 12.00 57.10 132.97 ;
        RECT 58.12 12.00 58.24 132.97 ;
        RECT 59.26 12.00 61.54 132.97 ;
        RECT 62.56 12.00 64.44 132.97 ;
        RECT 65.46 12.00 67.74 132.97 ;
        RECT 68.76 12.00 68.88 132.97 ;
        RECT 69.90 12.00 72.18 132.97 ;
        RECT 73.20 12.00 75.08 132.97 ;
        RECT 76.10 12.00 78.38 132.97 ;
        RECT 79.40 12.00 79.52 132.97 ;
        RECT 80.54 12.00 82.82 132.97 ;
        RECT 83.84 12.00 85.72 132.97 ;
        RECT 86.74 12.00 89.02 132.97 ;
        RECT 90.04 12.00 90.16 132.97 ;
        RECT 91.18 12.00 93.46 132.97 ;
        RECT 94.48 12.00 96.36 132.97 ;
        RECT 97.38 12.00 99.66 132.97 ;
        RECT 100.68 12.00 100.80 132.97 ;
        RECT 101.82 12.00 104.10 132.97 ;
        RECT 105.12 12.00 107.00 132.97 ;
        RECT 108.02 12.00 110.30 132.97 ;
        RECT 111.32 12.00 111.44 132.97 ;
        RECT 112.46 12.00 114.74 132.97 ;
        RECT 115.76 12.00 117.64 132.97 ;
        RECT 118.66 12.00 120.94 132.97 ;
        RECT 121.96 12.00 122.08 132.97 ;
        RECT 123.10 12.00 125.38 132.97 ;
        RECT 126.40 12.00 128.28 132.97 ;
        RECT 129.30 12.00 131.58 132.97 ;
        RECT 132.60 12.00 132.72 132.97 ;
        RECT 133.74 12.00 136.02 132.97 ;
        RECT 137.04 12.00 138.92 132.97 ;
        RECT 139.94 12.00 142.22 132.97 ;
        RECT 143.24 12.00 143.36 132.97 ;
        RECT 144.38 12.00 146.66 132.97 ;
        RECT 147.68 12.00 149.56 132.97 ;
        RECT 150.58 12.00 152.86 132.97 ;
        RECT 153.88 12.00 154.00 132.97 ;
        RECT 155.02 12.00 157.30 132.97 ;
        RECT 158.32 12.00 160.20 132.97 ;
        RECT 161.22 12.00 163.50 132.97 ;
        RECT 164.52 12.00 164.64 132.97 ;
        RECT 165.66 12.00 167.94 132.97 ;
        RECT 168.96 12.00 170.84 132.97 ;
        RECT 171.86 12.00 174.14 132.97 ;
        RECT 175.16 12.00 175.28 132.97 ;
        RECT 176.30 12.00 178.58 132.97 ;
        RECT 179.60 12.00 181.48 132.97 ;
        RECT 182.50 12.00 184.78 132.97 ;
        RECT 185.80 12.00 187.56 132.97 ;
        RECT 188.58 12.00 193.78 132.97 ;
        RECT 194.80 12.00 196.18 132.97 ;
        RECT 197.20 12.00 210.10 132.97 ;
        RECT 211.12 12.00 212.50 132.97 ;
        RECT 213.52 12.00 218.73 132.97 ;
        RECT 219.74 12.00 221.50 132.97 ;
        RECT 222.52 12.00 224.80 132.97 ;
        RECT 225.82 12.00 227.70 132.97 ;
        RECT 228.72 12.00 231.00 132.97 ;
        RECT 232.02 12.00 232.14 132.97 ;
        RECT 233.16 12.00 235.44 132.97 ;
        RECT 236.46 12.00 238.34 132.97 ;
        RECT 239.36 12.00 241.64 132.97 ;
        RECT 242.66 12.00 242.78 132.97 ;
        RECT 243.80 12.00 246.08 132.97 ;
        RECT 247.10 12.00 248.98 132.97 ;
        RECT 250.00 12.00 252.28 132.97 ;
        RECT 253.30 12.00 253.42 132.97 ;
        RECT 254.44 12.00 256.72 132.97 ;
        RECT 257.74 12.00 259.62 132.97 ;
        RECT 260.64 12.00 262.92 132.97 ;
        RECT 263.94 12.00 264.06 132.97 ;
        RECT 265.08 12.00 267.36 132.97 ;
        RECT 268.38 12.00 270.26 132.97 ;
        RECT 271.28 12.00 273.56 132.97 ;
        RECT 274.58 12.00 274.70 132.97 ;
        RECT 275.72 12.00 278.00 132.97 ;
        RECT 279.02 12.00 280.90 132.97 ;
        RECT 281.92 12.00 284.20 132.97 ;
        RECT 285.22 12.00 285.34 132.97 ;
        RECT 286.36 12.00 288.64 132.97 ;
        RECT 289.66 12.00 291.54 132.97 ;
        RECT 292.56 12.00 294.84 132.97 ;
        RECT 295.86 12.00 295.98 132.97 ;
        RECT 297.00 12.00 299.28 132.97 ;
        RECT 300.30 12.00 302.18 132.97 ;
        RECT 303.20 12.00 305.48 132.97 ;
        RECT 306.50 12.00 306.62 132.97 ;
        RECT 307.64 12.00 309.92 132.97 ;
        RECT 310.94 12.00 312.82 132.97 ;
        RECT 313.84 12.00 316.12 132.97 ;
        RECT 317.14 12.00 317.26 132.97 ;
        RECT 318.28 12.00 320.56 132.97 ;
        RECT 321.58 12.00 323.46 132.97 ;
        RECT 324.48 12.00 326.76 132.97 ;
        RECT 327.78 12.00 327.90 132.97 ;
        RECT 328.92 12.00 331.20 132.97 ;
        RECT 332.22 12.00 334.10 132.97 ;
        RECT 335.12 12.00 337.40 132.97 ;
        RECT 338.42 12.00 338.54 132.97 ;
        RECT 339.56 12.00 341.84 132.97 ;
        RECT 342.86 12.00 344.74 132.97 ;
        RECT 345.76 12.00 348.04 132.97 ;
        RECT 349.06 12.00 349.18 132.97 ;
        RECT 350.20 12.00 352.48 132.97 ;
        RECT 353.50 12.00 355.38 132.97 ;
        RECT 356.40 12.00 358.68 132.97 ;
        RECT 359.70 12.00 359.82 132.97 ;
        RECT 360.84 12.00 363.12 132.97 ;
        RECT 364.14 12.00 366.02 132.97 ;
        RECT 367.04 12.00 369.32 132.97 ;
        RECT 370.34 12.00 370.46 132.97 ;
        RECT 371.48 12.00 373.76 132.97 ;
        RECT 374.78 12.00 376.66 132.97 ;
        RECT 377.68 12.00 379.96 132.97 ;
        RECT 380.98 12.00 381.10 132.97 ;
        RECT 382.12 12.00 384.40 132.97 ;
        RECT 385.42 12.00 388.18 132.97 ;
        RECT 389.20 12.00 390.60 132.97 ;
        RECT 391.62 12.00 411.02 132.97 ;
        RECT 12.00 37.24 411.02 42.34 ;
        RECT 12.00 43.36 411.02 51.56 ;
        RECT 12.00 52.58 411.02 54.58 ;
        RECT 12.00 55.60 411.02 57.68 ;
        RECT 12.00 58.70 411.02 63.80 ;
        RECT 12.00 64.82 411.02 66.82 ;
        RECT 12.00 67.84 411.02 71.64 ;
        RECT 12.00 72.66 411.02 74.66 ;
        RECT 12.00 75.68 411.02 80.78 ;
        RECT 12.00 81.80 411.02 83.88 ;
        RECT 12.00 84.90 411.02 86.90 ;
        RECT 12.00 87.92 411.02 96.12 ;
        RECT 12.00 97.14 411.02 102.24 ;
        RECT 12.00 103.26 411.02 132.97 ;
    LAYER Metal4 ;
#      RECT 12.00 12.00 411.02 132.97 ;
        RECT 12.84 12.84 411.02 132.97 ;
        RECT 12.00 12.00 15.68 36.22 ;
        RECT 16.70 12.00 18.10 132.97 ;
        RECT 19.12 12.00 21.88 132.97 ;
        RECT 22.90 12.00 25.18 132.97 ;
        RECT 26.20 12.00 26.32 132.97 ;
        RECT 27.34 12.00 29.62 132.97 ;
        RECT 30.64 12.00 32.52 132.97 ;
        RECT 33.54 12.00 35.82 132.97 ;
        RECT 36.84 12.00 36.96 132.97 ;
        RECT 37.98 12.00 40.26 132.97 ;
        RECT 41.28 12.00 43.16 132.97 ;
        RECT 44.18 12.00 46.46 132.97 ;
        RECT 47.48 12.00 47.60 132.97 ;
        RECT 48.62 12.00 50.90 132.97 ;
        RECT 51.92 12.00 53.80 132.97 ;
        RECT 54.82 12.00 57.10 132.97 ;
        RECT 58.12 12.00 58.24 132.97 ;
        RECT 59.26 12.00 61.54 132.97 ;
        RECT 62.56 12.00 64.44 132.97 ;
        RECT 65.46 12.00 67.74 132.97 ;
        RECT 68.76 12.00 68.88 132.97 ;
        RECT 69.90 12.00 72.18 132.97 ;
        RECT 73.20 12.00 75.08 132.97 ;
        RECT 76.10 12.00 78.38 132.97 ;
        RECT 79.40 12.00 79.52 132.97 ;
        RECT 80.54 12.00 82.82 132.97 ;
        RECT 83.84 12.00 85.72 132.97 ;
        RECT 86.74 12.00 89.02 132.97 ;
        RECT 90.04 12.00 90.16 132.97 ;
        RECT 91.18 12.00 93.46 132.97 ;
        RECT 94.48 12.00 96.36 132.97 ;
        RECT 97.38 12.00 99.66 132.97 ;
        RECT 100.68 12.00 100.80 132.97 ;
        RECT 101.82 12.00 104.10 132.97 ;
        RECT 105.12 12.00 107.00 132.97 ;
        RECT 108.02 12.00 110.30 132.97 ;
        RECT 111.32 12.00 111.44 132.97 ;
        RECT 112.46 12.00 114.74 132.97 ;
        RECT 115.76 12.00 117.64 132.97 ;
        RECT 118.66 12.00 120.94 132.97 ;
        RECT 121.96 12.00 122.08 132.97 ;
        RECT 123.10 12.00 125.38 132.97 ;
        RECT 126.40 12.00 128.28 132.97 ;
        RECT 129.30 12.00 131.58 132.97 ;
        RECT 132.60 12.00 132.72 132.97 ;
        RECT 133.74 12.00 136.02 132.97 ;
        RECT 137.04 12.00 138.92 132.97 ;
        RECT 139.94 12.00 142.22 132.97 ;
        RECT 143.24 12.00 143.36 132.97 ;
        RECT 144.38 12.00 146.66 132.97 ;
        RECT 147.68 12.00 149.56 132.97 ;
        RECT 150.58 12.00 152.86 132.97 ;
        RECT 153.88 12.00 154.00 132.97 ;
        RECT 155.02 12.00 157.30 132.97 ;
        RECT 158.32 12.00 160.20 132.97 ;
        RECT 161.22 12.00 163.50 132.97 ;
        RECT 164.52 12.00 164.64 132.97 ;
        RECT 165.66 12.00 167.94 132.97 ;
        RECT 168.96 12.00 170.84 132.97 ;
        RECT 171.86 12.00 174.14 132.97 ;
        RECT 175.16 12.00 175.28 132.97 ;
        RECT 176.30 12.00 178.58 132.97 ;
        RECT 179.60 12.00 181.48 132.97 ;
        RECT 182.50 12.00 184.78 132.97 ;
        RECT 185.80 12.00 187.56 132.97 ;
        RECT 188.58 12.00 193.78 132.97 ;
        RECT 194.80 12.00 196.18 132.97 ;
        RECT 197.20 12.00 210.10 132.97 ;
        RECT 211.12 12.00 212.50 132.97 ;
        RECT 213.52 12.00 218.73 132.97 ;
        RECT 219.74 12.00 221.50 132.97 ;
        RECT 222.52 12.00 224.80 132.97 ;
        RECT 225.82 12.00 227.70 132.97 ;
        RECT 228.72 12.00 231.00 132.97 ;
        RECT 232.02 12.00 232.14 132.97 ;
        RECT 233.16 12.00 235.44 132.97 ;
        RECT 236.46 12.00 238.34 132.97 ;
        RECT 239.36 12.00 241.64 132.97 ;
        RECT 242.66 12.00 242.78 132.97 ;
        RECT 243.80 12.00 246.08 132.97 ;
        RECT 247.10 12.00 248.98 132.97 ;
        RECT 250.00 12.00 252.28 132.97 ;
        RECT 253.30 12.00 253.42 132.97 ;
        RECT 254.44 12.00 256.72 132.97 ;
        RECT 257.74 12.00 259.62 132.97 ;
        RECT 260.64 12.00 262.92 132.97 ;
        RECT 263.94 12.00 264.06 132.97 ;
        RECT 265.08 12.00 267.36 132.97 ;
        RECT 268.38 12.00 270.26 132.97 ;
        RECT 271.28 12.00 273.56 132.97 ;
        RECT 274.58 12.00 274.70 132.97 ;
        RECT 275.72 12.00 278.00 132.97 ;
        RECT 279.02 12.00 280.90 132.97 ;
        RECT 281.92 12.00 284.20 132.97 ;
        RECT 285.22 12.00 285.34 132.97 ;
        RECT 286.36 12.00 288.64 132.97 ;
        RECT 289.66 12.00 291.54 132.97 ;
        RECT 292.56 12.00 294.84 132.97 ;
        RECT 295.86 12.00 295.98 132.97 ;
        RECT 297.00 12.00 299.28 132.97 ;
        RECT 300.30 12.00 302.18 132.97 ;
        RECT 303.20 12.00 305.48 132.97 ;
        RECT 306.50 12.00 306.62 132.97 ;
        RECT 307.64 12.00 309.92 132.97 ;
        RECT 310.94 12.00 312.82 132.97 ;
        RECT 313.84 12.00 316.12 132.97 ;
        RECT 317.14 12.00 317.26 132.97 ;
        RECT 318.28 12.00 320.56 132.97 ;
        RECT 321.58 12.00 323.46 132.97 ;
        RECT 324.48 12.00 326.76 132.97 ;
        RECT 327.78 12.00 327.90 132.97 ;
        RECT 328.92 12.00 331.20 132.97 ;
        RECT 332.22 12.00 334.10 132.97 ;
        RECT 335.12 12.00 337.40 132.97 ;
        RECT 338.42 12.00 338.54 132.97 ;
        RECT 339.56 12.00 341.84 132.97 ;
        RECT 342.86 12.00 344.74 132.97 ;
        RECT 345.76 12.00 348.04 132.97 ;
        RECT 349.06 12.00 349.18 132.97 ;
        RECT 350.20 12.00 352.48 132.97 ;
        RECT 353.50 12.00 355.38 132.97 ;
        RECT 356.40 12.00 358.68 132.97 ;
        RECT 359.70 12.00 359.82 132.97 ;
        RECT 360.84 12.00 363.12 132.97 ;
        RECT 364.14 12.00 366.02 132.97 ;
        RECT 367.04 12.00 369.32 132.97 ;
        RECT 370.34 12.00 370.46 132.97 ;
        RECT 371.48 12.00 373.76 132.97 ;
        RECT 374.78 12.00 376.66 132.97 ;
        RECT 377.68 12.00 379.96 132.97 ;
        RECT 380.98 12.00 381.10 132.97 ;
        RECT 382.12 12.00 384.40 132.97 ;
        RECT 385.42 12.00 388.18 132.97 ;
        RECT 389.20 12.00 390.60 132.97 ;
        RECT 391.62 12.00 411.02 132.97 ;
        RECT 12.00 37.24 411.02 42.34 ;
        RECT 12.00 43.36 411.02 51.56 ;
        RECT 12.00 52.58 411.02 54.58 ;
        RECT 12.00 55.60 411.02 57.68 ;
        RECT 12.00 58.70 411.02 63.80 ;
        RECT 12.00 64.82 411.02 66.82 ;
        RECT 12.00 67.84 411.02 71.64 ;
        RECT 12.00 72.66 411.02 74.66 ;
        RECT 12.00 75.68 411.02 80.78 ;
        RECT 12.00 81.80 411.02 83.88 ;
        RECT 12.00 84.90 411.02 86.90 ;
        RECT 12.00 87.92 411.02 96.12 ;
        RECT 12.00 97.14 411.02 102.24 ;
        RECT 12.00 103.26 411.02 132.97 ;
    LAYER Metal5 ;
#      RECT 12.00 12.00 411.02 132.97 ;
        RECT 12.84 12.84 411.02 132.97 ;
        RECT 12.00 12.00 15.68 36.22 ;
        RECT 16.70 12.00 18.10 132.97 ;
        RECT 19.12 12.00 21.88 132.97 ;
        RECT 22.90 12.00 25.18 132.97 ;
        RECT 26.20 12.00 26.32 132.97 ;
        RECT 27.34 12.00 29.62 132.97 ;
        RECT 30.64 12.00 32.52 132.97 ;
        RECT 33.54 12.00 35.82 132.97 ;
        RECT 36.84 12.00 36.96 132.97 ;
        RECT 37.98 12.00 40.26 132.97 ;
        RECT 41.28 12.00 43.16 132.97 ;
        RECT 44.18 12.00 46.46 132.97 ;
        RECT 47.48 12.00 47.60 132.97 ;
        RECT 48.62 12.00 50.90 132.97 ;
        RECT 51.92 12.00 53.80 132.97 ;
        RECT 54.82 12.00 57.10 132.97 ;
        RECT 58.12 12.00 58.24 132.97 ;
        RECT 59.26 12.00 61.54 132.97 ;
        RECT 62.56 12.00 64.44 132.97 ;
        RECT 65.46 12.00 67.74 132.97 ;
        RECT 68.76 12.00 68.88 132.97 ;
        RECT 69.90 12.00 72.18 132.97 ;
        RECT 73.20 12.00 75.08 132.97 ;
        RECT 76.10 12.00 78.38 132.97 ;
        RECT 79.40 12.00 79.52 132.97 ;
        RECT 80.54 12.00 82.82 132.97 ;
        RECT 83.84 12.00 85.72 132.97 ;
        RECT 86.74 12.00 89.02 132.97 ;
        RECT 90.04 12.00 90.16 132.97 ;
        RECT 91.18 12.00 93.46 132.97 ;
        RECT 94.48 12.00 96.36 132.97 ;
        RECT 97.38 12.00 99.66 132.97 ;
        RECT 100.68 12.00 100.80 132.97 ;
        RECT 101.82 12.00 104.10 132.97 ;
        RECT 105.12 12.00 107.00 132.97 ;
        RECT 108.02 12.00 110.30 132.97 ;
        RECT 111.32 12.00 111.44 132.97 ;
        RECT 112.46 12.00 114.74 132.97 ;
        RECT 115.76 12.00 117.64 132.97 ;
        RECT 118.66 12.00 120.94 132.97 ;
        RECT 121.96 12.00 122.08 132.97 ;
        RECT 123.10 12.00 125.38 132.97 ;
        RECT 126.40 12.00 128.28 132.97 ;
        RECT 129.30 12.00 131.58 132.97 ;
        RECT 132.60 12.00 132.72 132.97 ;
        RECT 133.74 12.00 136.02 132.97 ;
        RECT 137.04 12.00 138.92 132.97 ;
        RECT 139.94 12.00 142.22 132.97 ;
        RECT 143.24 12.00 143.36 132.97 ;
        RECT 144.38 12.00 146.66 132.97 ;
        RECT 147.68 12.00 149.56 132.97 ;
        RECT 150.58 12.00 152.86 132.97 ;
        RECT 153.88 12.00 154.00 132.97 ;
        RECT 155.02 12.00 157.30 132.97 ;
        RECT 158.32 12.00 160.20 132.97 ;
        RECT 161.22 12.00 163.50 132.97 ;
        RECT 164.52 12.00 164.64 132.97 ;
        RECT 165.66 12.00 167.94 132.97 ;
        RECT 168.96 12.00 170.84 132.97 ;
        RECT 171.86 12.00 174.14 132.97 ;
        RECT 175.16 12.00 175.28 132.97 ;
        RECT 176.30 12.00 178.58 132.97 ;
        RECT 179.60 12.00 181.48 132.97 ;
        RECT 182.50 12.00 184.78 132.97 ;
        RECT 185.80 12.00 187.56 132.97 ;
        RECT 188.58 12.00 193.78 132.97 ;
        RECT 194.80 12.00 196.18 132.97 ;
        RECT 197.20 12.00 210.10 132.97 ;
        RECT 211.12 12.00 212.50 132.97 ;
        RECT 213.52 12.00 218.73 132.97 ;
        RECT 219.74 12.00 221.50 132.97 ;
        RECT 222.52 12.00 224.80 132.97 ;
        RECT 225.82 12.00 227.70 132.97 ;
        RECT 228.72 12.00 231.00 132.97 ;
        RECT 232.02 12.00 232.14 132.97 ;
        RECT 233.16 12.00 235.44 132.97 ;
        RECT 236.46 12.00 238.34 132.97 ;
        RECT 239.36 12.00 241.64 132.97 ;
        RECT 242.66 12.00 242.78 132.97 ;
        RECT 243.80 12.00 246.08 132.97 ;
        RECT 247.10 12.00 248.98 132.97 ;
        RECT 250.00 12.00 252.28 132.97 ;
        RECT 253.30 12.00 253.42 132.97 ;
        RECT 254.44 12.00 256.72 132.97 ;
        RECT 257.74 12.00 259.62 132.97 ;
        RECT 260.64 12.00 262.92 132.97 ;
        RECT 263.94 12.00 264.06 132.97 ;
        RECT 265.08 12.00 267.36 132.97 ;
        RECT 268.38 12.00 270.26 132.97 ;
        RECT 271.28 12.00 273.56 132.97 ;
        RECT 274.58 12.00 274.70 132.97 ;
        RECT 275.72 12.00 278.00 132.97 ;
        RECT 279.02 12.00 280.90 132.97 ;
        RECT 281.92 12.00 284.20 132.97 ;
        RECT 285.22 12.00 285.34 132.97 ;
        RECT 286.36 12.00 288.64 132.97 ;
        RECT 289.66 12.00 291.54 132.97 ;
        RECT 292.56 12.00 294.84 132.97 ;
        RECT 295.86 12.00 295.98 132.97 ;
        RECT 297.00 12.00 299.28 132.97 ;
        RECT 300.30 12.00 302.18 132.97 ;
        RECT 303.20 12.00 305.48 132.97 ;
        RECT 306.50 12.00 306.62 132.97 ;
        RECT 307.64 12.00 309.92 132.97 ;
        RECT 310.94 12.00 312.82 132.97 ;
        RECT 313.84 12.00 316.12 132.97 ;
        RECT 317.14 12.00 317.26 132.97 ;
        RECT 318.28 12.00 320.56 132.97 ;
        RECT 321.58 12.00 323.46 132.97 ;
        RECT 324.48 12.00 326.76 132.97 ;
        RECT 327.78 12.00 327.90 132.97 ;
        RECT 328.92 12.00 331.20 132.97 ;
        RECT 332.22 12.00 334.10 132.97 ;
        RECT 335.12 12.00 337.40 132.97 ;
        RECT 338.42 12.00 338.54 132.97 ;
        RECT 339.56 12.00 341.84 132.97 ;
        RECT 342.86 12.00 344.74 132.97 ;
        RECT 345.76 12.00 348.04 132.97 ;
        RECT 349.06 12.00 349.18 132.97 ;
        RECT 350.20 12.00 352.48 132.97 ;
        RECT 353.50 12.00 355.38 132.97 ;
        RECT 356.40 12.00 358.68 132.97 ;
        RECT 359.70 12.00 359.82 132.97 ;
        RECT 360.84 12.00 363.12 132.97 ;
        RECT 364.14 12.00 366.02 132.97 ;
        RECT 367.04 12.00 369.32 132.97 ;
        RECT 370.34 12.00 370.46 132.97 ;
        RECT 371.48 12.00 373.76 132.97 ;
        RECT 374.78 12.00 376.66 132.97 ;
        RECT 377.68 12.00 379.96 132.97 ;
        RECT 380.98 12.00 381.10 132.97 ;
        RECT 382.12 12.00 384.40 132.97 ;
        RECT 385.42 12.00 388.18 132.97 ;
        RECT 389.20 12.00 390.60 132.97 ;
        RECT 391.62 12.00 411.02 132.97 ;
        RECT 12.00 37.24 411.02 42.34 ;
        RECT 12.00 43.36 411.02 51.56 ;
        RECT 12.00 52.58 411.02 54.58 ;
        RECT 12.00 55.60 411.02 57.68 ;
        RECT 12.00 58.70 411.02 63.80 ;
        RECT 12.00 64.82 411.02 66.82 ;
        RECT 12.00 67.84 411.02 71.64 ;
        RECT 12.00 72.66 411.02 74.66 ;
        RECT 12.00 75.68 411.02 80.78 ;
        RECT 12.00 81.80 411.02 83.88 ;
        RECT 12.00 84.90 411.02 86.90 ;
        RECT 12.00 87.92 411.02 96.12 ;
        RECT 12.00 97.14 411.02 102.24 ;
        RECT 12.00 103.26 411.02 132.97 ;
    LAYER Metal6 ;
#      RECT 12.00 12.00 411.02 132.97 ;
        RECT 12.84 12.84 411.02 132.97 ;
        RECT 12.00 12.00 15.68 36.22 ;
        RECT 16.70 12.00 18.10 132.97 ;
        RECT 19.12 12.00 21.88 132.97 ;
        RECT 22.90 12.00 25.18 132.97 ;
        RECT 26.20 12.00 26.32 132.97 ;
        RECT 27.34 12.00 29.62 132.97 ;
        RECT 30.64 12.00 32.52 132.97 ;
        RECT 33.54 12.00 35.82 132.97 ;
        RECT 36.84 12.00 36.96 132.97 ;
        RECT 37.98 12.00 40.26 132.97 ;
        RECT 41.28 12.00 43.16 132.97 ;
        RECT 44.18 12.00 46.46 132.97 ;
        RECT 47.48 12.00 47.60 132.97 ;
        RECT 48.62 12.00 50.90 132.97 ;
        RECT 51.92 12.00 53.80 132.97 ;
        RECT 54.82 12.00 57.10 132.97 ;
        RECT 58.12 12.00 58.24 132.97 ;
        RECT 59.26 12.00 61.54 132.97 ;
        RECT 62.56 12.00 64.44 132.97 ;
        RECT 65.46 12.00 67.74 132.97 ;
        RECT 68.76 12.00 68.88 132.97 ;
        RECT 69.90 12.00 72.18 132.97 ;
        RECT 73.20 12.00 75.08 132.97 ;
        RECT 76.10 12.00 78.38 132.97 ;
        RECT 79.40 12.00 79.52 132.97 ;
        RECT 80.54 12.00 82.82 132.97 ;
        RECT 83.84 12.00 85.72 132.97 ;
        RECT 86.74 12.00 89.02 132.97 ;
        RECT 90.04 12.00 90.16 132.97 ;
        RECT 91.18 12.00 93.46 132.97 ;
        RECT 94.48 12.00 96.36 132.97 ;
        RECT 97.38 12.00 99.66 132.97 ;
        RECT 100.68 12.00 100.80 132.97 ;
        RECT 101.82 12.00 104.10 132.97 ;
        RECT 105.12 12.00 107.00 132.97 ;
        RECT 108.02 12.00 110.30 132.97 ;
        RECT 111.32 12.00 111.44 132.97 ;
        RECT 112.46 12.00 114.74 132.97 ;
        RECT 115.76 12.00 117.64 132.97 ;
        RECT 118.66 12.00 120.94 132.97 ;
        RECT 121.96 12.00 122.08 132.97 ;
        RECT 123.10 12.00 125.38 132.97 ;
        RECT 126.40 12.00 128.28 132.97 ;
        RECT 129.30 12.00 131.58 132.97 ;
        RECT 132.60 12.00 132.72 132.97 ;
        RECT 133.74 12.00 136.02 132.97 ;
        RECT 137.04 12.00 138.92 132.97 ;
        RECT 139.94 12.00 142.22 132.97 ;
        RECT 143.24 12.00 143.36 132.97 ;
        RECT 144.38 12.00 146.66 132.97 ;
        RECT 147.68 12.00 149.56 132.97 ;
        RECT 150.58 12.00 152.86 132.97 ;
        RECT 153.88 12.00 154.00 132.97 ;
        RECT 155.02 12.00 157.30 132.97 ;
        RECT 158.32 12.00 160.20 132.97 ;
        RECT 161.22 12.00 163.50 132.97 ;
        RECT 164.52 12.00 164.64 132.97 ;
        RECT 165.66 12.00 167.94 132.97 ;
        RECT 168.96 12.00 170.84 132.97 ;
        RECT 171.86 12.00 174.14 132.97 ;
        RECT 175.16 12.00 175.28 132.97 ;
        RECT 176.30 12.00 178.58 132.97 ;
        RECT 179.60 12.00 181.48 132.97 ;
        RECT 182.50 12.00 184.78 132.97 ;
        RECT 185.80 12.00 187.56 132.97 ;
        RECT 188.58 12.00 193.78 132.97 ;
        RECT 194.80 12.00 196.18 132.97 ;
        RECT 197.20 12.00 210.10 132.97 ;
        RECT 211.12 12.00 212.50 132.97 ;
        RECT 213.52 12.00 218.73 132.97 ;
        RECT 219.74 12.00 221.50 132.97 ;
        RECT 222.52 12.00 224.80 132.97 ;
        RECT 225.82 12.00 227.70 132.97 ;
        RECT 228.72 12.00 231.00 132.97 ;
        RECT 232.02 12.00 232.14 132.97 ;
        RECT 233.16 12.00 235.44 132.97 ;
        RECT 236.46 12.00 238.34 132.97 ;
        RECT 239.36 12.00 241.64 132.97 ;
        RECT 242.66 12.00 242.78 132.97 ;
        RECT 243.80 12.00 246.08 132.97 ;
        RECT 247.10 12.00 248.98 132.97 ;
        RECT 250.00 12.00 252.28 132.97 ;
        RECT 253.30 12.00 253.42 132.97 ;
        RECT 254.44 12.00 256.72 132.97 ;
        RECT 257.74 12.00 259.62 132.97 ;
        RECT 260.64 12.00 262.92 132.97 ;
        RECT 263.94 12.00 264.06 132.97 ;
        RECT 265.08 12.00 267.36 132.97 ;
        RECT 268.38 12.00 270.26 132.97 ;
        RECT 271.28 12.00 273.56 132.97 ;
        RECT 274.58 12.00 274.70 132.97 ;
        RECT 275.72 12.00 278.00 132.97 ;
        RECT 279.02 12.00 280.90 132.97 ;
        RECT 281.92 12.00 284.20 132.97 ;
        RECT 285.22 12.00 285.34 132.97 ;
        RECT 286.36 12.00 288.64 132.97 ;
        RECT 289.66 12.00 291.54 132.97 ;
        RECT 292.56 12.00 294.84 132.97 ;
        RECT 295.86 12.00 295.98 132.97 ;
        RECT 297.00 12.00 299.28 132.97 ;
        RECT 300.30 12.00 302.18 132.97 ;
        RECT 303.20 12.00 305.48 132.97 ;
        RECT 306.50 12.00 306.62 132.97 ;
        RECT 307.64 12.00 309.92 132.97 ;
        RECT 310.94 12.00 312.82 132.97 ;
        RECT 313.84 12.00 316.12 132.97 ;
        RECT 317.14 12.00 317.26 132.97 ;
        RECT 318.28 12.00 320.56 132.97 ;
        RECT 321.58 12.00 323.46 132.97 ;
        RECT 324.48 12.00 326.76 132.97 ;
        RECT 327.78 12.00 327.90 132.97 ;
        RECT 328.92 12.00 331.20 132.97 ;
        RECT 332.22 12.00 334.10 132.97 ;
        RECT 335.12 12.00 337.40 132.97 ;
        RECT 338.42 12.00 338.54 132.97 ;
        RECT 339.56 12.00 341.84 132.97 ;
        RECT 342.86 12.00 344.74 132.97 ;
        RECT 345.76 12.00 348.04 132.97 ;
        RECT 349.06 12.00 349.18 132.97 ;
        RECT 350.20 12.00 352.48 132.97 ;
        RECT 353.50 12.00 355.38 132.97 ;
        RECT 356.40 12.00 358.68 132.97 ;
        RECT 359.70 12.00 359.82 132.97 ;
        RECT 360.84 12.00 363.12 132.97 ;
        RECT 364.14 12.00 366.02 132.97 ;
        RECT 367.04 12.00 369.32 132.97 ;
        RECT 370.34 12.00 370.46 132.97 ;
        RECT 371.48 12.00 373.76 132.97 ;
        RECT 374.78 12.00 376.66 132.97 ;
        RECT 377.68 12.00 379.96 132.97 ;
        RECT 380.98 12.00 381.10 132.97 ;
        RECT 382.12 12.00 384.40 132.97 ;
        RECT 385.42 12.00 388.18 132.97 ;
        RECT 389.20 12.00 390.60 132.97 ;
        RECT 391.62 12.00 411.02 132.97 ;
        RECT 12.00 37.24 411.02 42.34 ;
        RECT 12.00 43.36 411.02 51.56 ;
        RECT 12.00 52.58 411.02 54.58 ;
        RECT 12.00 55.60 411.02 57.68 ;
        RECT 12.00 58.70 411.02 63.80 ;
        RECT 12.00 64.82 411.02 66.82 ;
        RECT 12.00 67.84 411.02 71.64 ;
        RECT 12.00 72.66 411.02 74.66 ;
        RECT 12.00 75.68 411.02 80.78 ;
        RECT 12.00 81.80 411.02 83.88 ;
        RECT 12.00 84.90 411.02 86.90 ;
        RECT 12.00 87.92 411.02 96.12 ;
        RECT 12.00 97.14 411.02 102.24 ;
        RECT 12.00 103.26 411.02 132.97 ;
  END
END MEM2


END LIBRARY

